module CPU6502Core(
  input         clock,
  input         reset,
  output [15:0] io_memAddr,
  output [7:0]  io_memDataOut,
  input  [7:0]  io_memDataIn,
  output        io_memWrite,
  output        io_memRead,
  output [7:0]  io_debug_regA,
  output [7:0]  io_debug_regX,
  output [7:0]  io_debug_regY,
  output [15:0] io_debug_regPC,
  output [7:0]  io_debug_regSP,
  output        io_debug_flagC,
  output        io_debug_flagZ,
  output        io_debug_flagN,
  output        io_debug_flagV,
  output [7:0]  io_debug_opcode
);
  reg [7:0] regs_a; // @[CPU6502Core.scala 19:21]
  reg [7:0] regs_x; // @[CPU6502Core.scala 19:21]
  reg [7:0] regs_y; // @[CPU6502Core.scala 19:21]
  reg [7:0] regs_sp; // @[CPU6502Core.scala 19:21]
  reg [15:0] regs_pc; // @[CPU6502Core.scala 19:21]
  reg  regs_flagC; // @[CPU6502Core.scala 19:21]
  reg  regs_flagZ; // @[CPU6502Core.scala 19:21]
  reg  regs_flagI; // @[CPU6502Core.scala 19:21]
  reg  regs_flagD; // @[CPU6502Core.scala 19:21]
  reg  regs_flagV; // @[CPU6502Core.scala 19:21]
  reg  regs_flagN; // @[CPU6502Core.scala 19:21]
  reg [1:0] state; // @[CPU6502Core.scala 23:22]
  reg [7:0] opcode; // @[CPU6502Core.scala 25:24]
  reg [15:0] operand; // @[CPU6502Core.scala 26:24]
  reg [2:0] cycle; // @[CPU6502Core.scala 27:24]
  wire [15:0] _regs_pc_T_1 = regs_pc + 16'h1; // @[CPU6502Core.scala 45:26]
  wire  _execResult_T = 8'h18 == opcode; // @[CPU6502Core.scala 89:20]
  wire  _execResult_T_1 = 8'h38 == opcode; // @[CPU6502Core.scala 89:20]
  wire  _execResult_T_2 = 8'hd8 == opcode; // @[CPU6502Core.scala 89:20]
  wire  _execResult_T_3 = 8'hf8 == opcode; // @[CPU6502Core.scala 89:20]
  wire  _execResult_T_4 = 8'h58 == opcode; // @[CPU6502Core.scala 89:20]
  wire  _execResult_T_5 = 8'h78 == opcode; // @[CPU6502Core.scala 89:20]
  wire  _execResult_T_6 = 8'hb8 == opcode; // @[CPU6502Core.scala 89:20]
  wire  _GEN_0 = _execResult_T_6 ? 1'h0 : regs_flagV; // @[Flag.scala 14:13 24:20 31:34]
  wire  _GEN_1 = _execResult_T_5 | regs_flagI; // @[Flag.scala 14:13 24:20 30:34]
  wire  _GEN_2 = _execResult_T_5 ? regs_flagV : _GEN_0; // @[Flag.scala 14:13 24:20]
  wire  _GEN_3 = _execResult_T_4 ? 1'h0 : _GEN_1; // @[Flag.scala 24:20 29:34]
  wire  _GEN_4 = _execResult_T_4 ? regs_flagV : _GEN_2; // @[Flag.scala 14:13 24:20]
  wire  _GEN_5 = _execResult_T_3 | regs_flagD; // @[Flag.scala 14:13 24:20 28:34]
  wire  _GEN_6 = _execResult_T_3 ? regs_flagI : _GEN_3; // @[Flag.scala 14:13 24:20]
  wire  _GEN_7 = _execResult_T_3 ? regs_flagV : _GEN_4; // @[Flag.scala 14:13 24:20]
  wire  _GEN_8 = _execResult_T_2 ? 1'h0 : _GEN_5; // @[Flag.scala 24:20 27:34]
  wire  _GEN_9 = _execResult_T_2 ? regs_flagI : _GEN_6; // @[Flag.scala 14:13 24:20]
  wire  _GEN_10 = _execResult_T_2 ? regs_flagV : _GEN_7; // @[Flag.scala 14:13 24:20]
  wire  _GEN_11 = _execResult_T_1 | regs_flagC; // @[Flag.scala 14:13 24:20 26:34]
  wire  _GEN_12 = _execResult_T_1 ? regs_flagD : _GEN_8; // @[Flag.scala 14:13 24:20]
  wire  _GEN_13 = _execResult_T_1 ? regs_flagI : _GEN_9; // @[Flag.scala 14:13 24:20]
  wire  _GEN_14 = _execResult_T_1 ? regs_flagV : _GEN_10; // @[Flag.scala 14:13 24:20]
  wire  execResult_result_newRegs_flagC = _execResult_T ? 1'h0 : _GEN_11; // @[Flag.scala 24:20 25:34]
  wire  execResult_result_newRegs_flagD = _execResult_T ? regs_flagD : _GEN_12; // @[Flag.scala 14:13 24:20]
  wire  execResult_result_newRegs_flagI = _execResult_T ? regs_flagI : _GEN_13; // @[Flag.scala 14:13 24:20]
  wire  execResult_result_newRegs_flagV = _execResult_T ? regs_flagV : _GEN_14; // @[Flag.scala 14:13 24:20]
  wire  _execResult_T_15 = 8'haa == opcode; // @[CPU6502Core.scala 89:20]
  wire  _execResult_T_16 = 8'ha8 == opcode; // @[CPU6502Core.scala 89:20]
  wire  _execResult_T_17 = 8'h8a == opcode; // @[CPU6502Core.scala 89:20]
  wire  _execResult_T_18 = 8'h98 == opcode; // @[CPU6502Core.scala 89:20]
  wire  _execResult_T_19 = 8'hba == opcode; // @[CPU6502Core.scala 89:20]
  wire  _execResult_T_20 = 8'h9a == opcode; // @[CPU6502Core.scala 89:20]
  wire  _execResult_result_newRegs_flagZ_T = regs_a == 8'h0; // @[Transfer.scala 28:33]
  wire [7:0] _GEN_19 = _execResult_T_20 ? regs_x : regs_sp; // @[Transfer.scala 14:13 24:20 51:20]
  wire [7:0] _GEN_20 = _execResult_T_19 ? regs_sp : regs_x; // @[Transfer.scala 14:13 24:20 46:19]
  wire  _GEN_21 = _execResult_T_19 ? regs_sp[7] : regs_flagN; // @[Transfer.scala 14:13 24:20 47:23]
  wire  _GEN_22 = _execResult_T_19 ? regs_sp == 8'h0 : regs_flagZ; // @[Transfer.scala 14:13 24:20 48:23]
  wire [7:0] _GEN_23 = _execResult_T_19 ? regs_sp : _GEN_19; // @[Transfer.scala 14:13 24:20]
  wire [7:0] _GEN_24 = _execResult_T_18 ? regs_y : regs_a; // @[Transfer.scala 14:13 24:20 41:19]
  wire  _GEN_25 = _execResult_T_18 ? regs_y[7] : _GEN_21; // @[Transfer.scala 24:20 42:23]
  wire  _GEN_26 = _execResult_T_18 ? regs_y == 8'h0 : _GEN_22; // @[Transfer.scala 24:20 43:23]
  wire [7:0] _GEN_27 = _execResult_T_18 ? regs_x : _GEN_20; // @[Transfer.scala 14:13 24:20]
  wire [7:0] _GEN_28 = _execResult_T_18 ? regs_sp : _GEN_23; // @[Transfer.scala 14:13 24:20]
  wire [7:0] _GEN_29 = _execResult_T_17 ? regs_x : _GEN_24; // @[Transfer.scala 24:20 36:19]
  wire  _GEN_30 = _execResult_T_17 ? regs_x[7] : _GEN_25; // @[Transfer.scala 24:20 37:23]
  wire  _GEN_31 = _execResult_T_17 ? regs_x == 8'h0 : _GEN_26; // @[Transfer.scala 24:20 38:23]
  wire [7:0] _GEN_32 = _execResult_T_17 ? regs_x : _GEN_27; // @[Transfer.scala 14:13 24:20]
  wire [7:0] _GEN_33 = _execResult_T_17 ? regs_sp : _GEN_28; // @[Transfer.scala 14:13 24:20]
  wire [7:0] _GEN_34 = _execResult_T_16 ? regs_a : regs_y; // @[Transfer.scala 14:13 24:20 31:19]
  wire  _GEN_35 = _execResult_T_16 ? regs_a[7] : _GEN_30; // @[Transfer.scala 24:20 32:23]
  wire  _GEN_36 = _execResult_T_16 ? _execResult_result_newRegs_flagZ_T : _GEN_31; // @[Transfer.scala 24:20 33:23]
  wire [7:0] _GEN_37 = _execResult_T_16 ? regs_a : _GEN_29; // @[Transfer.scala 14:13 24:20]
  wire [7:0] _GEN_38 = _execResult_T_16 ? regs_x : _GEN_32; // @[Transfer.scala 14:13 24:20]
  wire [7:0] _GEN_39 = _execResult_T_16 ? regs_sp : _GEN_33; // @[Transfer.scala 14:13 24:20]
  wire [7:0] execResult_result_newRegs_1_x = _execResult_T_15 ? regs_a : _GEN_38; // @[Transfer.scala 24:20 26:19]
  wire  execResult_result_newRegs_1_flagN = _execResult_T_15 ? regs_a[7] : _GEN_35; // @[Transfer.scala 24:20 27:23]
  wire  execResult_result_newRegs_1_flagZ = _execResult_T_15 ? regs_a == 8'h0 : _GEN_36; // @[Transfer.scala 24:20 28:23]
  wire [7:0] execResult_result_newRegs_1_y = _execResult_T_15 ? regs_y : _GEN_34; // @[Transfer.scala 14:13 24:20]
  wire [7:0] execResult_result_newRegs_1_a = _execResult_T_15 ? regs_a : _GEN_37; // @[Transfer.scala 14:13 24:20]
  wire [7:0] execResult_result_newRegs_1_sp = _execResult_T_15 ? regs_sp : _GEN_39; // @[Transfer.scala 14:13 24:20]
  wire  _execResult_T_26 = 8'he8 == opcode; // @[CPU6502Core.scala 89:20]
  wire  _execResult_T_27 = 8'hc8 == opcode; // @[CPU6502Core.scala 89:20]
  wire  _execResult_T_28 = 8'hca == opcode; // @[CPU6502Core.scala 89:20]
  wire  _execResult_T_29 = 8'h88 == opcode; // @[CPU6502Core.scala 89:20]
  wire  _execResult_T_30 = 8'h1a == opcode; // @[CPU6502Core.scala 89:20]
  wire  _execResult_T_31 = 8'h3a == opcode; // @[CPU6502Core.scala 89:20]
  wire [7:0] execResult_result_res = regs_x + 8'h1; // @[Arithmetic.scala 34:26]
  wire [7:0] execResult_result_res_1 = regs_y + 8'h1; // @[Arithmetic.scala 40:26]
  wire [7:0] execResult_result_res_2 = regs_x - 8'h1; // @[Arithmetic.scala 46:26]
  wire [7:0] execResult_result_res_3 = regs_y - 8'h1; // @[Arithmetic.scala 52:26]
  wire [7:0] execResult_result_res_4 = regs_a + 8'h1; // @[Arithmetic.scala 58:26]
  wire [7:0] execResult_result_res_5 = regs_a - 8'h1; // @[Arithmetic.scala 64:26]
  wire [7:0] _GEN_46 = _execResult_T_31 ? execResult_result_res_5 : regs_a; // @[Arithmetic.scala 22:13 32:20 65:19]
  wire  _GEN_47 = _execResult_T_31 ? execResult_result_res_5[7] : regs_flagN; // @[Arithmetic.scala 22:13 32:20 66:23]
  wire  _GEN_48 = _execResult_T_31 ? execResult_result_res_5 == 8'h0 : regs_flagZ; // @[Arithmetic.scala 22:13 32:20 67:23]
  wire [7:0] _GEN_49 = _execResult_T_30 ? execResult_result_res_4 : _GEN_46; // @[Arithmetic.scala 32:20 59:19]
  wire  _GEN_50 = _execResult_T_30 ? execResult_result_res_4[7] : _GEN_47; // @[Arithmetic.scala 32:20 60:23]
  wire  _GEN_51 = _execResult_T_30 ? execResult_result_res_4 == 8'h0 : _GEN_48; // @[Arithmetic.scala 32:20 61:23]
  wire [7:0] _GEN_52 = _execResult_T_29 ? execResult_result_res_3 : regs_y; // @[Arithmetic.scala 22:13 32:20 53:19]
  wire  _GEN_53 = _execResult_T_29 ? execResult_result_res_3[7] : _GEN_50; // @[Arithmetic.scala 32:20 54:23]
  wire  _GEN_54 = _execResult_T_29 ? execResult_result_res_3 == 8'h0 : _GEN_51; // @[Arithmetic.scala 32:20 55:23]
  wire [7:0] _GEN_55 = _execResult_T_29 ? regs_a : _GEN_49; // @[Arithmetic.scala 22:13 32:20]
  wire [7:0] _GEN_56 = _execResult_T_28 ? execResult_result_res_2 : regs_x; // @[Arithmetic.scala 22:13 32:20 47:19]
  wire  _GEN_57 = _execResult_T_28 ? execResult_result_res_2[7] : _GEN_53; // @[Arithmetic.scala 32:20 48:23]
  wire  _GEN_58 = _execResult_T_28 ? execResult_result_res_2 == 8'h0 : _GEN_54; // @[Arithmetic.scala 32:20 49:23]
  wire [7:0] _GEN_59 = _execResult_T_28 ? regs_y : _GEN_52; // @[Arithmetic.scala 22:13 32:20]
  wire [7:0] _GEN_60 = _execResult_T_28 ? regs_a : _GEN_55; // @[Arithmetic.scala 22:13 32:20]
  wire [7:0] _GEN_61 = _execResult_T_27 ? execResult_result_res_1 : _GEN_59; // @[Arithmetic.scala 32:20 41:19]
  wire  _GEN_62 = _execResult_T_27 ? execResult_result_res_1[7] : _GEN_57; // @[Arithmetic.scala 32:20 42:23]
  wire  _GEN_63 = _execResult_T_27 ? execResult_result_res_1 == 8'h0 : _GEN_58; // @[Arithmetic.scala 32:20 43:23]
  wire [7:0] _GEN_64 = _execResult_T_27 ? regs_x : _GEN_56; // @[Arithmetic.scala 22:13 32:20]
  wire [7:0] _GEN_65 = _execResult_T_27 ? regs_a : _GEN_60; // @[Arithmetic.scala 22:13 32:20]
  wire [7:0] execResult_result_newRegs_2_x = _execResult_T_26 ? execResult_result_res : _GEN_64; // @[Arithmetic.scala 32:20 35:19]
  wire  execResult_result_newRegs_2_flagN = _execResult_T_26 ? execResult_result_res[7] : _GEN_62; // @[Arithmetic.scala 32:20 36:23]
  wire  execResult_result_newRegs_2_flagZ = _execResult_T_26 ? execResult_result_res == 8'h0 : _GEN_63; // @[Arithmetic.scala 32:20 37:23]
  wire [7:0] execResult_result_newRegs_2_y = _execResult_T_26 ? regs_y : _GEN_61; // @[Arithmetic.scala 22:13 32:20]
  wire [7:0] execResult_result_newRegs_2_a = _execResult_T_26 ? regs_a : _GEN_65; // @[Arithmetic.scala 22:13 32:20]
  wire [8:0] _execResult_result_sum_T = regs_a + io_memDataIn; // @[Arithmetic.scala 81:22]
  wire [8:0] _GEN_1508 = {{8'd0}, regs_flagC}; // @[Arithmetic.scala 81:35]
  wire [9:0] execResult_result_sum = _execResult_result_sum_T + _GEN_1508; // @[Arithmetic.scala 81:35]
  wire [7:0] execResult_result_newRegs_3_a = execResult_result_sum[7:0]; // @[Arithmetic.scala 82:21]
  wire  execResult_result_newRegs_3_flagC = execResult_result_sum[8]; // @[Arithmetic.scala 83:25]
  wire  execResult_result_newRegs_3_flagN = execResult_result_sum[7]; // @[Arithmetic.scala 84:25]
  wire  execResult_result_newRegs_3_flagZ = execResult_result_newRegs_3_a == 8'h0; // @[Arithmetic.scala 85:32]
  wire  execResult_result_newRegs_3_flagV = regs_a[7] == io_memDataIn[7] & regs_a[7] !=
    execResult_result_newRegs_3_flagN; // @[Arithmetic.scala 86:51]
  wire [8:0] _execResult_result_diff_T = regs_a - io_memDataIn; // @[Arithmetic.scala 106:23]
  wire  _execResult_result_diff_T_2 = ~regs_flagC; // @[Arithmetic.scala 106:40]
  wire [8:0] _GEN_1509 = {{8'd0}, _execResult_result_diff_T_2}; // @[Arithmetic.scala 106:36]
  wire [9:0] execResult_result_diff = _execResult_result_diff_T - _GEN_1509; // @[Arithmetic.scala 106:36]
  wire [7:0] execResult_result_newRegs_4_a = execResult_result_diff[7:0]; // @[Arithmetic.scala 107:22]
  wire  execResult_result_newRegs_4_flagC = ~execResult_result_diff[8]; // @[Arithmetic.scala 108:22]
  wire  execResult_result_newRegs_4_flagN = execResult_result_diff[7]; // @[Arithmetic.scala 109:26]
  wire  execResult_result_newRegs_4_flagZ = execResult_result_newRegs_4_a == 8'h0; // @[Arithmetic.scala 110:33]
  wire  execResult_result_newRegs_4_flagV = regs_a[7] != io_memDataIn[7] & regs_a[7] !=
    execResult_result_newRegs_4_flagN; // @[Arithmetic.scala 111:51]
  wire [2:0] _execResult_result_result_nextCycle_T_1 = cycle + 3'h1; // @[Arithmetic.scala 132:31]
  wire  _execResult_result_T_20 = 3'h0 == cycle; // @[Arithmetic.scala 140:19]
  wire  _execResult_result_T_21 = 3'h1 == cycle; // @[Arithmetic.scala 140:19]
  wire  _execResult_result_T_22 = 3'h2 == cycle; // @[Arithmetic.scala 140:19]
  wire [7:0] _execResult_result_res_T_8 = io_memDataIn + 8'h1; // @[Arithmetic.scala 156:52]
  wire [7:0] _execResult_result_res_T_10 = io_memDataIn - 8'h1; // @[Arithmetic.scala 156:69]
  wire [7:0] execResult_result_res_6 = opcode == 8'he6 ? _execResult_result_res_T_8 : _execResult_result_res_T_10; // @[Arithmetic.scala 156:22]
  wire [15:0] _GEN_71 = 3'h2 == cycle ? operand : 16'h0; // @[Arithmetic.scala 140:19 134:20 155:24]
  wire [7:0] _GEN_72 = 3'h2 == cycle ? execResult_result_res_6 : 8'h0; // @[Arithmetic.scala 140:19 135:20 157:24]
  wire  _GEN_74 = 3'h2 == cycle ? execResult_result_res_6[7] : regs_flagN; // @[Arithmetic.scala 129:13 140:19 159:23]
  wire  _GEN_75 = 3'h2 == cycle ? execResult_result_res_6 == 8'h0 : regs_flagZ; // @[Arithmetic.scala 129:13 140:19 160:23]
  wire [15:0] execResult_result_newRegs_5_pc = 3'h0 == cycle ? _regs_pc_T_1 : regs_pc; // @[Arithmetic.scala 129:13 140:19 145:20]
  wire  _GEN_94 = 3'h1 == cycle ? regs_flagZ : _GEN_75; // @[Arithmetic.scala 129:13 140:19]
  wire  execResult_result_newRegs_5_flagZ = 3'h0 == cycle ? regs_flagZ : _GEN_94; // @[Arithmetic.scala 129:13 140:19]
  wire  _GEN_93 = 3'h1 == cycle ? regs_flagN : _GEN_74; // @[Arithmetic.scala 129:13 140:19]
  wire  execResult_result_newRegs_5_flagN = 3'h0 == cycle ? regs_flagN : _GEN_93; // @[Arithmetic.scala 129:13 140:19]
  wire [15:0] _GEN_88 = 3'h1 == cycle ? operand : _GEN_71; // @[Arithmetic.scala 140:19 150:24]
  wire [2:0] _GEN_90 = 3'h1 == cycle ? 3'h2 : _execResult_result_result_nextCycle_T_1; // @[Arithmetic.scala 140:19 132:22 152:26]
  wire [7:0] _GEN_91 = 3'h1 == cycle ? 8'h0 : _GEN_72; // @[Arithmetic.scala 140:19 135:20]
  wire  _GEN_92 = 3'h1 == cycle ? 1'h0 : 3'h2 == cycle; // @[Arithmetic.scala 140:19 136:21]
  wire [15:0] execResult_result_result_6_memAddr = 3'h0 == cycle ? regs_pc : _GEN_88; // @[Arithmetic.scala 140:19 142:24]
  wire  execResult_result_result_6_memRead = 3'h0 == cycle | 3'h1 == cycle; // @[Arithmetic.scala 140:19 143:24]
  wire [15:0] execResult_result_result_6_operand = 3'h0 == cycle ? {{8'd0}, io_memDataIn} : operand; // @[Arithmetic.scala 140:19 138:20 144:24]
  wire [2:0] execResult_result_result_6_nextCycle = 3'h0 == cycle ? 3'h1 : _GEN_90; // @[Arithmetic.scala 140:19 147:26]
  wire [7:0] execResult_result_result_6_memData = 3'h0 == cycle ? 8'h0 : _GEN_91; // @[Arithmetic.scala 140:19 135:20]
  wire  execResult_result_result_6_done = 3'h0 == cycle ? 1'h0 : _GEN_92; // @[Arithmetic.scala 140:19 136:21]
  wire  _execResult_T_42 = 8'h29 == opcode; // @[CPU6502Core.scala 89:20]
  wire  _execResult_T_43 = 8'h9 == opcode; // @[CPU6502Core.scala 89:20]
  wire  _execResult_T_44 = 8'h49 == opcode; // @[CPU6502Core.scala 89:20]
  wire [7:0] _execResult_result_res_T_11 = regs_a & io_memDataIn; // @[Logic.scala 24:34]
  wire [7:0] _execResult_result_res_T_12 = regs_a | io_memDataIn; // @[Logic.scala 25:34]
  wire [7:0] _execResult_result_res_T_13 = regs_a ^ io_memDataIn; // @[Logic.scala 26:34]
  wire [7:0] _GEN_128 = _execResult_T_44 ? _execResult_result_res_T_13 : 8'h0; // @[Logic.scala 23:20 26:24 21:9]
  wire [7:0] _GEN_129 = _execResult_T_43 ? _execResult_result_res_T_12 : _GEN_128; // @[Logic.scala 23:20 25:24]
  wire [7:0] execResult_result_res_7 = _execResult_T_42 ? _execResult_result_res_T_11 : _GEN_129; // @[Logic.scala 23:20 24:24]
  wire  execResult_result_newRegs_6_flagN = execResult_result_res_7[7]; // @[Logic.scala 30:25]
  wire  execResult_result_newRegs_6_flagZ = execResult_result_res_7 == 8'h0; // @[Logic.scala 31:26]
  wire [15:0] _GEN_131 = _execResult_result_T_21 ? operand : 16'h0; // @[Logic.scala 60:19 54:20 70:24]
  wire  _GEN_133 = _execResult_result_T_21 ? _execResult_result_res_T_11 == 8'h0 : regs_flagZ; // @[Logic.scala 49:13 60:19 72:23]
  wire  _GEN_134 = _execResult_result_T_21 ? io_memDataIn[7] : regs_flagN; // @[Logic.scala 49:13 60:19 73:23]
  wire  _GEN_135 = _execResult_result_T_21 ? io_memDataIn[6] : regs_flagV; // @[Logic.scala 49:13 60:19 74:23]
  wire  execResult_result_newRegs_7_flagZ = _execResult_result_T_20 ? regs_flagZ : _GEN_133; // @[Logic.scala 49:13 60:19]
  wire  execResult_result_newRegs_7_flagV = _execResult_result_T_20 ? regs_flagV : _GEN_135; // @[Logic.scala 49:13 60:19]
  wire  execResult_result_newRegs_7_flagN = _execResult_result_T_20 ? regs_flagN : _GEN_134; // @[Logic.scala 49:13 60:19]
  wire [15:0] execResult_result_result_8_memAddr = _execResult_result_T_20 ? regs_pc : _GEN_131; // @[Logic.scala 60:19 62:24]
  wire [2:0] execResult_result_result_8_nextCycle = _execResult_result_T_20 ? 3'h1 :
    _execResult_result_result_nextCycle_T_1; // @[Logic.scala 60:19 52:22 67:26]
  wire  execResult_result_result_8_done = _execResult_result_T_20 ? 1'h0 : _execResult_result_T_21; // @[Logic.scala 51:17 60:19]
  wire  _execResult_T_48 = 8'ha == opcode; // @[CPU6502Core.scala 89:20]
  wire  _execResult_T_49 = 8'h4a == opcode; // @[CPU6502Core.scala 89:20]
  wire  _execResult_T_50 = 8'h2a == opcode; // @[CPU6502Core.scala 89:20]
  wire  _execResult_T_51 = 8'h6a == opcode; // @[CPU6502Core.scala 89:20]
  wire [8:0] _execResult_result_res_T_14 = {regs_a, 1'h0}; // @[Shift.scala 35:24]
  wire [7:0] _execResult_result_res_T_18 = {regs_a[6:0],regs_flagC}; // @[Cat.scala 33:92]
  wire [7:0] _execResult_result_res_T_20 = {regs_flagC,regs_a[7:1]}; // @[Cat.scala 33:92]
  wire  _GEN_169 = _execResult_T_51 ? regs_a[0] : regs_flagC; // @[Shift.scala 18:13 32:20 46:23]
  wire [7:0] _GEN_170 = _execResult_T_51 ? _execResult_result_res_T_20 : regs_a; // @[Shift.scala 32:20 47:13 29:9]
  wire  _GEN_171 = _execResult_T_50 ? regs_a[7] : _GEN_169; // @[Shift.scala 32:20 42:23]
  wire [7:0] _GEN_172 = _execResult_T_50 ? _execResult_result_res_T_18 : _GEN_170; // @[Shift.scala 32:20 43:13]
  wire  _GEN_173 = _execResult_T_49 ? regs_a[0] : _GEN_171; // @[Shift.scala 32:20 38:23]
  wire [7:0] _GEN_174 = _execResult_T_49 ? {{1'd0}, regs_a[7:1]} : _GEN_172; // @[Shift.scala 32:20 39:13]
  wire  execResult_result_newRegs_8_flagC = _execResult_T_48 ? regs_a[7] : _GEN_173; // @[Shift.scala 32:20 34:23]
  wire [7:0] execResult_result_res_8 = _execResult_T_48 ? _execResult_result_res_T_14[7:0] : _GEN_174; // @[Shift.scala 32:20 35:13]
  wire  execResult_result_newRegs_8_flagN = execResult_result_res_8[7]; // @[Shift.scala 52:25]
  wire  execResult_result_newRegs_8_flagZ = execResult_result_res_8 == 8'h0; // @[Shift.scala 53:26]
  wire  _execResult_T_55 = 8'h6 == opcode; // @[CPU6502Core.scala 89:20]
  wire  _execResult_T_56 = 8'h46 == opcode; // @[CPU6502Core.scala 89:20]
  wire  _execResult_T_57 = 8'h26 == opcode; // @[CPU6502Core.scala 89:20]
  wire  _execResult_T_58 = 8'h66 == opcode; // @[CPU6502Core.scala 89:20]
  wire [8:0] _execResult_result_res_T_21 = {io_memDataIn, 1'h0}; // @[Shift.scala 95:31]
  wire [7:0] _execResult_result_res_T_25 = {io_memDataIn[6:0],regs_flagC}; // @[Cat.scala 33:92]
  wire [7:0] _execResult_result_res_T_27 = {regs_flagC,io_memDataIn[7:1]}; // @[Cat.scala 33:92]
  wire  _GEN_177 = _execResult_T_58 ? io_memDataIn[0] : regs_flagC; // @[Shift.scala 92:24 108:27 62:13]
  wire [7:0] _GEN_178 = _execResult_T_58 ? _execResult_result_res_T_27 : 8'h0; // @[Shift.scala 109:17 90:13 92:24]
  wire  _GEN_179 = _execResult_T_57 ? io_memDataIn[7] : _GEN_177; // @[Shift.scala 92:24 103:27]
  wire [7:0] _GEN_180 = _execResult_T_57 ? _execResult_result_res_T_25 : _GEN_178; // @[Shift.scala 104:17 92:24]
  wire  _GEN_181 = _execResult_T_56 ? io_memDataIn[0] : _GEN_179; // @[Shift.scala 92:24 98:27]
  wire [7:0] _GEN_182 = _execResult_T_56 ? {{1'd0}, io_memDataIn[7:1]} : _GEN_180; // @[Shift.scala 92:24 99:17]
  wire  _GEN_183 = _execResult_T_55 ? io_memDataIn[7] : _GEN_181; // @[Shift.scala 92:24 94:27]
  wire [7:0] execResult_result_res_9 = _execResult_T_55 ? _execResult_result_res_T_21[7:0] : _GEN_182; // @[Shift.scala 92:24 95:17]
  wire  _GEN_186 = _execResult_result_T_22 ? _GEN_183 : regs_flagC; // @[Shift.scala 62:13 73:19]
  wire [7:0] _GEN_187 = _execResult_result_T_22 ? execResult_result_res_9 : 8'h0; // @[Shift.scala 73:19 113:24 68:20]
  wire  _GEN_189 = _execResult_result_T_22 ? execResult_result_res_9[7] : regs_flagN; // @[Shift.scala 73:19 115:23 62:13]
  wire  _GEN_190 = _execResult_result_T_22 ? execResult_result_res_9 == 8'h0 : regs_flagZ; // @[Shift.scala 73:19 116:23 62:13]
  wire  _GEN_206 = _execResult_result_T_21 ? regs_flagC : _GEN_186; // @[Shift.scala 62:13 73:19]
  wire  execResult_result_newRegs_9_flagC = _execResult_result_T_20 ? regs_flagC : _GEN_206; // @[Shift.scala 62:13 73:19]
  wire  _GEN_210 = _execResult_result_T_21 ? regs_flagZ : _GEN_190; // @[Shift.scala 62:13 73:19]
  wire  execResult_result_newRegs_9_flagZ = _execResult_result_T_20 ? regs_flagZ : _GEN_210; // @[Shift.scala 62:13 73:19]
  wire  _GEN_209 = _execResult_result_T_21 ? regs_flagN : _GEN_189; // @[Shift.scala 62:13 73:19]
  wire  execResult_result_newRegs_9_flagN = _execResult_result_T_20 ? regs_flagN : _GEN_209; // @[Shift.scala 62:13 73:19]
  wire [7:0] _GEN_207 = _execResult_result_T_21 ? 8'h0 : _GEN_187; // @[Shift.scala 73:19 68:20]
  wire [7:0] execResult_result_result_10_memData = _execResult_result_T_20 ? 8'h0 : _GEN_207; // @[Shift.scala 73:19 68:20]
  wire  _execResult_T_62 = 8'hc9 == opcode; // @[CPU6502Core.scala 89:20]
  wire  _execResult_T_63 = 8'he0 == opcode; // @[CPU6502Core.scala 89:20]
  wire  _execResult_T_64 = 8'hc0 == opcode; // @[CPU6502Core.scala 89:20]
  wire [7:0] _GEN_245 = _execResult_T_64 ? regs_y : regs_a; // @[Compare.scala 21:14 23:20 26:29]
  wire [7:0] _GEN_246 = _execResult_T_63 ? regs_x : _GEN_245; // @[Compare.scala 23:20 25:29]
  wire [7:0] execResult_result_regValue = _execResult_T_62 ? regs_a : _GEN_246; // @[Compare.scala 23:20 24:29]
  wire [8:0] execResult_result_diff_1 = execResult_result_regValue - io_memDataIn; // @[Compare.scala 29:25]
  wire  execResult_result_newRegs_10_flagC = execResult_result_regValue >= io_memDataIn; // @[Compare.scala 30:31]
  wire  execResult_result_newRegs_10_flagZ = execResult_result_regValue == io_memDataIn; // @[Compare.scala 31:31]
  wire  execResult_result_newRegs_10_flagN = execResult_result_diff_1[7]; // @[Compare.scala 32:26]
  wire  _GEN_250 = _execResult_result_T_21 ? regs_a >= io_memDataIn : regs_flagC; // @[Compare.scala 50:13 61:19 74:23]
  wire  _GEN_251 = _execResult_result_T_21 ? regs_a == io_memDataIn : regs_flagZ; // @[Compare.scala 50:13 61:19 75:23]
  wire  _GEN_252 = _execResult_result_T_21 ? _execResult_result_diff_T[7] : regs_flagN; // @[Compare.scala 50:13 61:19 76:23]
  wire  execResult_result_newRegs_11_flagC = _execResult_result_T_20 ? regs_flagC : _GEN_250; // @[Compare.scala 50:13 61:19]
  wire  execResult_result_newRegs_11_flagZ = _execResult_result_T_20 ? regs_flagZ : _GEN_251; // @[Compare.scala 50:13 61:19]
  wire  execResult_result_newRegs_11_flagN = _execResult_result_T_20 ? regs_flagN : _GEN_252; // @[Compare.scala 50:13 61:19]
  wire  _execResult_T_68 = 8'hf0 == opcode; // @[CPU6502Core.scala 89:20]
  wire  _execResult_T_69 = 8'hd0 == opcode; // @[CPU6502Core.scala 89:20]
  wire  _execResult_T_70 = 8'hb0 == opcode; // @[CPU6502Core.scala 89:20]
  wire  _execResult_T_71 = 8'h90 == opcode; // @[CPU6502Core.scala 89:20]
  wire  _execResult_T_72 = 8'h30 == opcode; // @[CPU6502Core.scala 89:20]
  wire  _execResult_T_73 = 8'h10 == opcode; // @[CPU6502Core.scala 89:20]
  wire  _execResult_T_74 = 8'h50 == opcode; // @[CPU6502Core.scala 89:20]
  wire  _execResult_T_75 = 8'h70 == opcode; // @[CPU6502Core.scala 89:20]
  wire  _GEN_286 = _execResult_T_74 & ~regs_flagV; // @[Branch.scala 18:16 20:20 28:31]
  wire  _GEN_287 = _execResult_T_75 ? regs_flagV : _GEN_286; // @[Branch.scala 20:20 27:31]
  wire  _GEN_288 = _execResult_T_73 ? ~regs_flagN : _GEN_287; // @[Branch.scala 20:20 26:31]
  wire  _GEN_289 = _execResult_T_72 ? regs_flagN : _GEN_288; // @[Branch.scala 20:20 25:31]
  wire  _GEN_290 = _execResult_T_71 ? _execResult_result_diff_T_2 : _GEN_289; // @[Branch.scala 20:20 24:31]
  wire  _GEN_291 = _execResult_T_70 ? regs_flagC : _GEN_290; // @[Branch.scala 20:20 23:31]
  wire  _GEN_292 = _execResult_T_69 ? ~regs_flagZ : _GEN_291; // @[Branch.scala 20:20 22:31]
  wire  execResult_result_takeBranch = _execResult_T_68 ? regs_flagZ : _GEN_292; // @[Branch.scala 20:20 21:31]
  wire [7:0] execResult_result_offset = io_memDataIn; // @[Branch.scala 32:28]
  wire [15:0] _execResult_result_newRegs_pc_T_16 = regs_pc + 16'h1; // @[Branch.scala 34:43]
  wire [15:0] _GEN_1510 = {{8{execResult_result_offset[7]}},execResult_result_offset}; // @[Branch.scala 34:50]
  wire [15:0] _execResult_result_newRegs_pc_T_20 = $signed(_execResult_result_newRegs_pc_T_16) + $signed(_GEN_1510); // @[Branch.scala 34:60]
  wire [15:0] execResult_result_newRegs_12_pc = execResult_result_takeBranch ? _execResult_result_newRegs_pc_T_20 :
    _regs_pc_T_1; // @[Branch.scala 34:22]
  wire  _execResult_T_83 = 8'ha9 == opcode; // @[CPU6502Core.scala 89:20]
  wire  _execResult_T_84 = 8'ha2 == opcode; // @[CPU6502Core.scala 89:20]
  wire  _execResult_T_85 = 8'ha0 == opcode; // @[CPU6502Core.scala 89:20]
  wire [7:0] _GEN_294 = _execResult_T_85 ? io_memDataIn : regs_y; // @[LoadStore.scala 23:13 25:20 28:30]
  wire [7:0] _GEN_295 = _execResult_T_84 ? io_memDataIn : regs_x; // @[LoadStore.scala 23:13 25:20 27:30]
  wire [7:0] _GEN_296 = _execResult_T_84 ? regs_y : _GEN_294; // @[LoadStore.scala 23:13 25:20]
  wire [7:0] execResult_result_newRegs_13_a = _execResult_T_83 ? io_memDataIn : regs_a; // @[LoadStore.scala 23:13 25:20 26:30]
  wire [7:0] execResult_result_newRegs_13_x = _execResult_T_83 ? regs_x : _GEN_295; // @[LoadStore.scala 23:13 25:20]
  wire [7:0] execResult_result_newRegs_13_y = _execResult_T_83 ? regs_y : _GEN_296; // @[LoadStore.scala 23:13 25:20]
  wire  execResult_result_newRegs_13_flagZ = io_memDataIn == 8'h0; // @[LoadStore.scala 32:32]
  wire  execResult_result_isLoad = opcode == 8'ha5; // @[LoadStore.scala 61:25]
  wire  execResult_result_isStoreA = opcode == 8'h85; // @[LoadStore.scala 62:27]
  wire  execResult_result_isStoreX = opcode == 8'h86; // @[LoadStore.scala 63:27]
  wire [7:0] _execResult_result_result_memData_T = execResult_result_isStoreX ? regs_x : regs_y; // @[LoadStore.scala 84:54]
  wire [7:0] _execResult_result_result_memData_T_1 = execResult_result_isStoreA ? regs_a :
    _execResult_result_result_memData_T; // @[LoadStore.scala 84:32]
  wire [7:0] _GEN_301 = execResult_result_isLoad ? io_memDataIn : regs_a; // @[LoadStore.scala 50:13 77:22 79:21]
  wire  _GEN_302 = execResult_result_isLoad ? io_memDataIn[7] : regs_flagN; // @[LoadStore.scala 50:13 77:22 80:25]
  wire  _GEN_303 = execResult_result_isLoad ? execResult_result_newRegs_13_flagZ : regs_flagZ; // @[LoadStore.scala 50:13 77:22 81:25]
  wire  _GEN_304 = execResult_result_isLoad ? 1'h0 : 1'h1; // @[LoadStore.scala 57:21 77:22 83:27]
  wire [7:0] _GEN_305 = execResult_result_isLoad ? 8'h0 : _execResult_result_result_memData_T_1; // @[LoadStore.scala 56:20 77:22 84:26]
  wire  _GEN_307 = _execResult_result_T_21 & execResult_result_isLoad; // @[LoadStore.scala 66:19 58:20]
  wire [7:0] _GEN_308 = _execResult_result_T_21 ? _GEN_301 : regs_a; // @[LoadStore.scala 50:13 66:19]
  wire  _GEN_309 = _execResult_result_T_21 ? _GEN_302 : regs_flagN; // @[LoadStore.scala 50:13 66:19]
  wire  _GEN_310 = _execResult_result_T_21 ? _GEN_303 : regs_flagZ; // @[LoadStore.scala 50:13 66:19]
  wire [7:0] _GEN_312 = _execResult_result_T_21 ? _GEN_305 : 8'h0; // @[LoadStore.scala 66:19 56:20]
  wire [7:0] execResult_result_newRegs_14_a = _execResult_result_T_20 ? regs_a : _GEN_308; // @[LoadStore.scala 50:13 66:19]
  wire  execResult_result_newRegs_14_flagZ = _execResult_result_T_20 ? regs_flagZ : _GEN_310; // @[LoadStore.scala 50:13 66:19]
  wire  execResult_result_newRegs_14_flagN = _execResult_result_T_20 ? regs_flagN : _GEN_309; // @[LoadStore.scala 50:13 66:19]
  wire  execResult_result_result_15_memRead = _execResult_result_T_20 | _GEN_307; // @[LoadStore.scala 66:19 69:24]
  wire  execResult_result_result_15_memWrite = _execResult_result_T_20 ? 1'h0 : _execResult_result_T_21 & _GEN_304; // @[LoadStore.scala 66:19 57:21]
  wire [7:0] execResult_result_result_15_memData = _execResult_result_T_20 ? 8'h0 : _GEN_312; // @[LoadStore.scala 66:19 56:20]
  wire  execResult_result_isLoad_1 = opcode == 8'hb5; // @[LoadStore.scala 109:25]
  wire [7:0] _execResult_result_result_operand_T_1 = io_memDataIn + regs_x; // @[LoadStore.scala 115:38]
  wire [7:0] _GEN_350 = execResult_result_isLoad_1 ? io_memDataIn : regs_a; // @[LoadStore.scala 122:22 124:21 98:13]
  wire  _GEN_351 = execResult_result_isLoad_1 ? io_memDataIn[7] : regs_flagN; // @[LoadStore.scala 122:22 125:25 98:13]
  wire  _GEN_352 = execResult_result_isLoad_1 ? execResult_result_newRegs_13_flagZ : regs_flagZ; // @[LoadStore.scala 122:22 126:25 98:13]
  wire  _GEN_353 = execResult_result_isLoad_1 ? 1'h0 : 1'h1; // @[LoadStore.scala 105:21 122:22 128:27]
  wire [7:0] _GEN_354 = execResult_result_isLoad_1 ? 8'h0 : regs_a; // @[LoadStore.scala 104:20 122:22 129:26]
  wire  _GEN_356 = _execResult_result_T_21 & execResult_result_isLoad_1; // @[LoadStore.scala 111:19 106:20]
  wire [7:0] _GEN_357 = _execResult_result_T_21 ? _GEN_350 : regs_a; // @[LoadStore.scala 111:19 98:13]
  wire  _GEN_358 = _execResult_result_T_21 ? _GEN_351 : regs_flagN; // @[LoadStore.scala 111:19 98:13]
  wire  _GEN_359 = _execResult_result_T_21 ? _GEN_352 : regs_flagZ; // @[LoadStore.scala 111:19 98:13]
  wire [7:0] _GEN_361 = _execResult_result_T_21 ? _GEN_354 : 8'h0; // @[LoadStore.scala 111:19 104:20]
  wire [7:0] execResult_result_newRegs_15_a = _execResult_result_T_20 ? regs_a : _GEN_357; // @[LoadStore.scala 111:19 98:13]
  wire  execResult_result_newRegs_15_flagZ = _execResult_result_T_20 ? regs_flagZ : _GEN_359; // @[LoadStore.scala 111:19 98:13]
  wire  execResult_result_newRegs_15_flagN = _execResult_result_T_20 ? regs_flagN : _GEN_358; // @[LoadStore.scala 111:19 98:13]
  wire  execResult_result_result_16_memRead = _execResult_result_T_20 | _GEN_356; // @[LoadStore.scala 111:19 114:24]
  wire [15:0] execResult_result_result_16_operand = _execResult_result_T_20 ? {{8'd0},
    _execResult_result_result_operand_T_1} : operand; // @[LoadStore.scala 111:19 107:20 115:24]
  wire  execResult_result_result_16_memWrite = _execResult_result_T_20 ? 1'h0 : _execResult_result_T_21 & _GEN_353; // @[LoadStore.scala 111:19 105:21]
  wire [7:0] execResult_result_result_16_memData = _execResult_result_T_20 ? 8'h0 : _GEN_361; // @[LoadStore.scala 111:19 104:20]
  wire  execResult_result_isLoad_2 = opcode == 8'had; // @[LoadStore.scala 154:25]
  wire [15:0] _execResult_result_result_operand_T_4 = {io_memDataIn,operand[7:0]}; // @[Cat.scala 33:92]
  wire [7:0] _GEN_399 = execResult_result_isLoad_2 ? io_memDataIn : regs_a; // @[LoadStore.scala 143:13 175:22 177:21]
  wire  _GEN_400 = execResult_result_isLoad_2 ? io_memDataIn[7] : regs_flagN; // @[LoadStore.scala 143:13 175:22 178:25]
  wire  _GEN_401 = execResult_result_isLoad_2 ? execResult_result_newRegs_13_flagZ : regs_flagZ; // @[LoadStore.scala 143:13 175:22 179:25]
  wire  _GEN_402 = execResult_result_isLoad_2 ? 1'h0 : 1'h1; // @[LoadStore.scala 150:21 175:22 181:27]
  wire [7:0] _GEN_403 = execResult_result_isLoad_2 ? 8'h0 : regs_a; // @[LoadStore.scala 149:20 175:22 182:26]
  wire  _GEN_405 = _execResult_result_T_22 & execResult_result_isLoad_2; // @[LoadStore.scala 156:19 151:20]
  wire [7:0] _GEN_406 = _execResult_result_T_22 ? _GEN_399 : regs_a; // @[LoadStore.scala 143:13 156:19]
  wire  _GEN_407 = _execResult_result_T_22 ? _GEN_400 : regs_flagN; // @[LoadStore.scala 143:13 156:19]
  wire  _GEN_408 = _execResult_result_T_22 ? _GEN_401 : regs_flagZ; // @[LoadStore.scala 143:13 156:19]
  wire [7:0] _GEN_410 = _execResult_result_T_22 ? _GEN_403 : 8'h0; // @[LoadStore.scala 156:19 149:20]
  wire [7:0] _GEN_441 = _execResult_result_T_21 ? regs_a : _GEN_406; // @[LoadStore.scala 143:13 156:19]
  wire [7:0] execResult_result_newRegs_16_a = _execResult_result_T_20 ? regs_a : _GEN_441; // @[LoadStore.scala 143:13 156:19]
  wire [15:0] _GEN_427 = _execResult_result_T_21 ? _regs_pc_T_1 : regs_pc; // @[LoadStore.scala 143:13 156:19 169:20]
  wire [15:0] execResult_result_newRegs_16_pc = _execResult_result_T_20 ? _regs_pc_T_1 : _GEN_427; // @[LoadStore.scala 156:19 161:20]
  wire  _GEN_443 = _execResult_result_T_21 ? regs_flagZ : _GEN_408; // @[LoadStore.scala 143:13 156:19]
  wire  execResult_result_newRegs_16_flagZ = _execResult_result_T_20 ? regs_flagZ : _GEN_443; // @[LoadStore.scala 143:13 156:19]
  wire  _GEN_442 = _execResult_result_T_21 ? regs_flagN : _GEN_407; // @[LoadStore.scala 143:13 156:19]
  wire  execResult_result_newRegs_16_flagN = _execResult_result_T_20 ? regs_flagN : _GEN_442; // @[LoadStore.scala 143:13 156:19]
  wire [15:0] _GEN_424 = _execResult_result_T_21 ? regs_pc : _GEN_71; // @[LoadStore.scala 156:19 166:24]
  wire  _GEN_425 = _execResult_result_T_21 | _GEN_405; // @[LoadStore.scala 156:19 167:24]
  wire [15:0] _GEN_426 = _execResult_result_T_21 ? _execResult_result_result_operand_T_4 : operand; // @[LoadStore.scala 156:19 152:20 168:24]
  wire  _GEN_444 = _execResult_result_T_21 ? 1'h0 : _execResult_result_T_22 & _GEN_402; // @[LoadStore.scala 156:19 150:21]
  wire [7:0] _GEN_445 = _execResult_result_T_21 ? 8'h0 : _GEN_410; // @[LoadStore.scala 156:19 149:20]
  wire [15:0] execResult_result_result_17_memAddr = _execResult_result_T_20 ? regs_pc : _GEN_424; // @[LoadStore.scala 156:19 158:24]
  wire  execResult_result_result_17_memRead = _execResult_result_T_20 | _GEN_425; // @[LoadStore.scala 156:19 159:24]
  wire [15:0] execResult_result_result_17_operand = _execResult_result_T_20 ? {{8'd0}, io_memDataIn} : _GEN_426; // @[LoadStore.scala 156:19 160:24]
  wire  execResult_result_result_17_memWrite = _execResult_result_T_20 ? 1'h0 : _GEN_444; // @[LoadStore.scala 156:19 150:21]
  wire [7:0] execResult_result_result_17_memData = _execResult_result_T_20 ? 8'h0 : _GEN_445; // @[LoadStore.scala 156:19 149:20]
  wire [7:0] execResult_result_indexReg = opcode == 8'hbd ? regs_x : regs_y; // @[LoadStore.scala 207:23]
  wire [15:0] _GEN_1511 = {{8'd0}, execResult_result_indexReg}; // @[LoadStore.scala 221:57]
  wire [15:0] _execResult_result_result_operand_T_8 = _execResult_result_result_operand_T_4 + _GEN_1511; // @[LoadStore.scala 221:57]
  wire [7:0] _GEN_472 = _execResult_result_T_22 ? io_memDataIn : regs_a; // @[LoadStore.scala 196:13 209:19 229:19]
  wire  _GEN_473 = _execResult_result_T_22 ? io_memDataIn[7] : regs_flagN; // @[LoadStore.scala 196:13 209:19 230:23]
  wire  _GEN_474 = _execResult_result_T_22 ? execResult_result_newRegs_13_flagZ : regs_flagZ; // @[LoadStore.scala 196:13 209:19 231:23]
  wire [7:0] _GEN_504 = _execResult_result_T_21 ? regs_a : _GEN_472; // @[LoadStore.scala 196:13 209:19]
  wire [7:0] execResult_result_newRegs_17_a = _execResult_result_T_20 ? regs_a : _GEN_504; // @[LoadStore.scala 196:13 209:19]
  wire  _GEN_506 = _execResult_result_T_21 ? regs_flagZ : _GEN_474; // @[LoadStore.scala 196:13 209:19]
  wire  execResult_result_newRegs_17_flagZ = _execResult_result_T_20 ? regs_flagZ : _GEN_506; // @[LoadStore.scala 196:13 209:19]
  wire  _GEN_505 = _execResult_result_T_21 ? regs_flagN : _GEN_473; // @[LoadStore.scala 196:13 209:19]
  wire  execResult_result_newRegs_17_flagN = _execResult_result_T_20 ? regs_flagN : _GEN_505; // @[LoadStore.scala 196:13 209:19]
  wire  _GEN_488 = _execResult_result_T_21 | _execResult_result_T_22; // @[LoadStore.scala 209:19 220:24]
  wire [15:0] _GEN_489 = _execResult_result_T_21 ? _execResult_result_result_operand_T_8 : operand; // @[LoadStore.scala 209:19 205:20 221:24]
  wire  execResult_result_result_18_memRead = _execResult_result_T_20 | _GEN_488; // @[LoadStore.scala 209:19 212:24]
  wire [15:0] execResult_result_result_18_operand = _execResult_result_T_20 ? {{8'd0}, io_memDataIn} : _GEN_489; // @[LoadStore.scala 209:19 213:24]
  wire [7:0] _execResult_result_pushData_T = {regs_flagN,regs_flagV,2'h3,regs_flagD,regs_flagI,regs_flagZ,regs_flagC}; // @[Cat.scala 33:92]
  wire [7:0] execResult_result_pushData = opcode == 8'h8 ? _execResult_result_pushData_T : regs_a; // @[Stack.scala 21:14 23:29 24:16]
  wire [7:0] execResult_result_newRegs_18_sp = regs_sp - 8'h1; // @[Stack.scala 27:27]
  wire [15:0] execResult_result_result_19_memAddr = {8'h1,regs_sp}; // @[Cat.scala 33:92]
  wire [7:0] _execResult_result_newRegs_sp_T_3 = regs_sp + 8'h1; // @[Stack.scala 57:31]
  wire [7:0] _GEN_530 = opcode == 8'h68 ? io_memDataIn : regs_a; // @[Stack.scala 44:13 65:33 66:21]
  wire  _GEN_531 = opcode == 8'h68 ? io_memDataIn[7] : io_memDataIn[7]; // @[Stack.scala 65:33 67:25 75:25]
  wire  _GEN_532 = opcode == 8'h68 ? execResult_result_newRegs_13_flagZ : io_memDataIn[1]; // @[Stack.scala 65:33 68:25 71:25]
  wire  _GEN_533 = opcode == 8'h68 ? regs_flagC : io_memDataIn[0]; // @[Stack.scala 44:13 65:33 70:25]
  wire  _GEN_534 = opcode == 8'h68 ? regs_flagI : io_memDataIn[2]; // @[Stack.scala 44:13 65:33 72:25]
  wire  _GEN_535 = opcode == 8'h68 ? regs_flagD : io_memDataIn[3]; // @[Stack.scala 44:13 65:33 73:25]
  wire  _GEN_536 = opcode == 8'h68 ? regs_flagV : io_memDataIn[6]; // @[Stack.scala 44:13 65:33 74:25]
  wire [15:0] _GEN_537 = _execResult_result_T_21 ? execResult_result_result_19_memAddr : 16'h0; // @[Stack.scala 55:19 49:20 62:24]
  wire [7:0] _GEN_539 = _execResult_result_T_21 ? _GEN_530 : regs_a; // @[Stack.scala 44:13 55:19]
  wire  _GEN_540 = _execResult_result_T_21 ? _GEN_531 : regs_flagN; // @[Stack.scala 44:13 55:19]
  wire  _GEN_541 = _execResult_result_T_21 ? _GEN_532 : regs_flagZ; // @[Stack.scala 44:13 55:19]
  wire  _GEN_542 = _execResult_result_T_21 ? _GEN_533 : regs_flagC; // @[Stack.scala 44:13 55:19]
  wire  _GEN_543 = _execResult_result_T_21 ? _GEN_534 : regs_flagI; // @[Stack.scala 44:13 55:19]
  wire  _GEN_544 = _execResult_result_T_21 ? _GEN_535 : regs_flagD; // @[Stack.scala 44:13 55:19]
  wire  _GEN_545 = _execResult_result_T_21 ? _GEN_536 : regs_flagV; // @[Stack.scala 44:13 55:19]
  wire [7:0] execResult_result_newRegs_19_a = _execResult_result_T_20 ? regs_a : _GEN_539; // @[Stack.scala 44:13 55:19]
  wire [7:0] execResult_result_newRegs_19_sp = _execResult_result_T_20 ? _execResult_result_newRegs_sp_T_3 : regs_sp; // @[Stack.scala 44:13 55:19 57:20]
  wire  execResult_result_newRegs_19_flagC = _execResult_result_T_20 ? regs_flagC : _GEN_542; // @[Stack.scala 44:13 55:19]
  wire  execResult_result_newRegs_19_flagZ = _execResult_result_T_20 ? regs_flagZ : _GEN_541; // @[Stack.scala 44:13 55:19]
  wire  execResult_result_newRegs_19_flagI = _execResult_result_T_20 ? regs_flagI : _GEN_543; // @[Stack.scala 44:13 55:19]
  wire  execResult_result_newRegs_19_flagD = _execResult_result_T_20 ? regs_flagD : _GEN_544; // @[Stack.scala 44:13 55:19]
  wire  execResult_result_newRegs_19_flagV = _execResult_result_T_20 ? regs_flagV : _GEN_545; // @[Stack.scala 44:13 55:19]
  wire  execResult_result_newRegs_19_flagN = _execResult_result_T_20 ? regs_flagN : _GEN_540; // @[Stack.scala 44:13 55:19]
  wire [15:0] execResult_result_result_20_memAddr = _execResult_result_T_20 ? 16'h0 : _GEN_537; // @[Stack.scala 55:19 49:20]
  wire [15:0] _GEN_581 = _execResult_result_T_21 ? regs_pc : 16'h0; // @[Jump.scala 26:19 20:20 36:24]
  wire [15:0] _GEN_583 = _execResult_result_T_21 ? _execResult_result_result_operand_T_4 : regs_pc; // @[Jump.scala 15:13 26:19 38:20]
  wire [15:0] execResult_result_newRegs_20_pc = _execResult_result_T_20 ? _regs_pc_T_1 : _GEN_583; // @[Jump.scala 26:19 31:20]
  wire [15:0] execResult_result_result_21_memAddr = _execResult_result_T_20 ? regs_pc : _GEN_581; // @[Jump.scala 26:19 28:24]
  wire  _execResult_result_T_74 = 3'h3 == cycle; // @[Jump.scala 62:19]
  wire [15:0] _GEN_614 = 3'h3 == cycle ? execResult_result_result_19_memAddr : 16'h0; // @[Jump.scala 62:19 56:20 86:24]
  wire [7:0] _GEN_615 = 3'h3 == cycle ? regs_pc[7:0] : 8'h0; // @[Jump.scala 62:19 57:20 87:24]
  wire [7:0] _GEN_617 = 3'h3 == cycle ? execResult_result_newRegs_18_sp : regs_sp; // @[Jump.scala 51:13 62:19 89:20]
  wire [15:0] _GEN_618 = 3'h3 == cycle ? operand : regs_pc; // @[Jump.scala 51:13 62:19 90:20]
  wire [7:0] _GEN_634 = _execResult_result_T_22 ? execResult_result_newRegs_18_sp : _GEN_617; // @[Jump.scala 62:19 81:20]
  wire [7:0] _GEN_656 = _execResult_result_T_21 ? regs_sp : _GEN_634; // @[Jump.scala 51:13 62:19]
  wire [7:0] execResult_result_newRegs_21_sp = _execResult_result_T_20 ? regs_sp : _GEN_656; // @[Jump.scala 51:13 62:19]
  wire [15:0] _GEN_648 = _execResult_result_T_22 ? regs_pc : _GEN_618; // @[Jump.scala 51:13 62:19]
  wire [15:0] _GEN_669 = _execResult_result_T_21 ? regs_pc : _GEN_648; // @[Jump.scala 51:13 62:19]
  wire [15:0] execResult_result_newRegs_21_pc = _execResult_result_T_20 ? _regs_pc_T_1 : _GEN_669; // @[Jump.scala 62:19 67:20]
  wire [15:0] _GEN_631 = _execResult_result_T_22 ? execResult_result_result_19_memAddr : _GEN_614; // @[Jump.scala 62:19 78:24]
  wire [7:0] _GEN_632 = _execResult_result_T_22 ? regs_pc[15:8] : _GEN_615; // @[Jump.scala 62:19 79:24]
  wire  _GEN_633 = _execResult_result_T_22 | 3'h3 == cycle; // @[Jump.scala 62:19 80:25]
  wire [2:0] _GEN_647 = _execResult_result_T_22 ? 3'h3 : _execResult_result_result_nextCycle_T_1; // @[Jump.scala 62:19 54:22 83:26]
  wire  _GEN_649 = _execResult_result_T_22 ? 1'h0 : 3'h3 == cycle; // @[Jump.scala 53:17 62:19]
  wire [15:0] _GEN_650 = _execResult_result_T_21 ? regs_pc : _GEN_631; // @[Jump.scala 62:19 72:24]
  wire [2:0] _GEN_653 = _execResult_result_T_21 ? 3'h2 : _GEN_647; // @[Jump.scala 62:19 75:26]
  wire [7:0] _GEN_654 = _execResult_result_T_21 ? 8'h0 : _GEN_632; // @[Jump.scala 62:19 57:20]
  wire  _GEN_655 = _execResult_result_T_21 ? 1'h0 : _GEN_633; // @[Jump.scala 62:19 58:21]
  wire  _GEN_670 = _execResult_result_T_21 ? 1'h0 : _GEN_649; // @[Jump.scala 53:17 62:19]
  wire [15:0] execResult_result_result_22_memAddr = _execResult_result_T_20 ? regs_pc : _GEN_650; // @[Jump.scala 62:19 64:24]
  wire [2:0] execResult_result_result_22_nextCycle = _execResult_result_T_20 ? 3'h1 : _GEN_653; // @[Jump.scala 62:19 69:26]
  wire [7:0] execResult_result_result_22_memData = _execResult_result_T_20 ? 8'h0 : _GEN_654; // @[Jump.scala 62:19 57:20]
  wire  execResult_result_result_22_memWrite = _execResult_result_T_20 ? 1'h0 : _GEN_655; // @[Jump.scala 62:19 58:21]
  wire  execResult_result_result_22_done = _execResult_result_T_20 ? 1'h0 : _GEN_670; // @[Jump.scala 53:17 62:19]
  wire [15:0] _execResult_result_newRegs_pc_T_45 = _execResult_result_result_operand_T_4 + 16'h1; // @[Jump.scala 131:53]
  wire [15:0] _GEN_692 = _execResult_result_T_22 ? execResult_result_result_19_memAddr : 16'h0; // @[Jump.scala 114:19 108:20 129:24]
  wire [15:0] _GEN_694 = _execResult_result_T_22 ? _execResult_result_newRegs_pc_T_45 : regs_pc; // @[Jump.scala 103:13 114:19 131:20]
  wire [7:0] _GEN_710 = _execResult_result_T_21 ? _execResult_result_newRegs_sp_T_3 : regs_sp; // @[Jump.scala 103:13 114:19 124:20]
  wire [7:0] execResult_result_newRegs_22_sp = _execResult_result_T_20 ? _execResult_result_newRegs_sp_T_3 : _GEN_710; // @[Jump.scala 114:19 116:20]
  wire [15:0] _GEN_724 = _execResult_result_T_21 ? regs_pc : _GEN_694; // @[Jump.scala 103:13 114:19]
  wire [15:0] execResult_result_newRegs_22_pc = _execResult_result_T_20 ? regs_pc : _GEN_724; // @[Jump.scala 103:13 114:19]
  wire [15:0] _GEN_707 = _execResult_result_T_21 ? execResult_result_result_19_memAddr : _GEN_692; // @[Jump.scala 114:19 121:24]
  wire [15:0] _GEN_709 = _execResult_result_T_21 ? {{8'd0}, io_memDataIn} : operand; // @[Jump.scala 114:19 112:20 123:24]
  wire [15:0] execResult_result_result_23_memAddr = _execResult_result_T_20 ? 16'h0 : _GEN_707; // @[Jump.scala 114:19 108:20]
  wire  execResult_result_result_23_memRead = _execResult_result_T_20 ? 1'h0 : _GEN_488; // @[Jump.scala 114:19 111:20]
  wire [15:0] execResult_result_result_23_operand = _execResult_result_T_20 ? operand : _GEN_709; // @[Jump.scala 114:19 112:20]
  wire [15:0] _GEN_745 = 3'h5 == cycle ? 16'hffff : 16'h0; // @[Jump.scala 155:19 149:20 195:24]
  wire [15:0] _GEN_747 = 3'h5 == cycle ? _execResult_result_result_operand_T_4 : regs_pc; // @[Jump.scala 144:13 155:19 197:20]
  wire [7:0] _GEN_827 = _execResult_result_T_21 ? execResult_result_newRegs_18_sp : _GEN_634; // @[Jump.scala 155:19 165:20]
  wire [7:0] execResult_result_newRegs_23_sp = _execResult_result_T_20 ? regs_sp : _GEN_827; // @[Jump.scala 144:13 155:19]
  wire [15:0] _GEN_764 = 3'h4 == cycle ? regs_pc : _GEN_747; // @[Jump.scala 144:13 155:19]
  wire [15:0] _GEN_799 = _execResult_result_T_74 ? regs_pc : _GEN_764; // @[Jump.scala 144:13 155:19]
  wire [15:0] _GEN_822 = _execResult_result_T_22 ? regs_pc : _GEN_799; // @[Jump.scala 144:13 155:19]
  wire [15:0] _GEN_845 = _execResult_result_T_21 ? regs_pc : _GEN_822; // @[Jump.scala 144:13 155:19]
  wire [15:0] execResult_result_newRegs_23_pc = _execResult_result_T_20 ? _regs_pc_T_1 : _GEN_845; // @[Jump.scala 155:19 157:20]
  wire  _GEN_782 = _execResult_result_T_74 | regs_flagI; // @[Jump.scala 144:13 155:19 183:23]
  wire  _GEN_818 = _execResult_result_T_22 ? regs_flagI : _GEN_782; // @[Jump.scala 144:13 155:19]
  wire  _GEN_841 = _execResult_result_T_21 ? regs_flagI : _GEN_818; // @[Jump.scala 144:13 155:19]
  wire  execResult_result_newRegs_23_flagI = _execResult_result_T_20 ? regs_flagI : _GEN_841; // @[Jump.scala 144:13 155:19]
  wire [15:0] _GEN_760 = 3'h4 == cycle ? 16'hfffe : _GEN_745; // @[Jump.scala 155:19 189:24]
  wire  _GEN_761 = 3'h4 == cycle | 3'h5 == cycle; // @[Jump.scala 155:19 190:24]
  wire [15:0] _GEN_762 = 3'h4 == cycle ? {{8'd0}, io_memDataIn} : operand; // @[Jump.scala 155:19 153:20 191:24]
  wire [2:0] _GEN_763 = 3'h4 == cycle ? 3'h5 : _execResult_result_result_nextCycle_T_1; // @[Jump.scala 155:19 147:22 192:26]
  wire  _GEN_777 = 3'h4 == cycle ? 1'h0 : 3'h5 == cycle; // @[Jump.scala 146:17 155:19]
  wire [15:0] _GEN_778 = _execResult_result_T_74 ? execResult_result_result_19_memAddr : _GEN_760; // @[Jump.scala 155:19 179:24]
  wire [7:0] _GEN_779 = _execResult_result_T_74 ? _execResult_result_pushData_T : 8'h0; // @[Jump.scala 155:19 150:20 180:24]
  wire [2:0] _GEN_796 = _execResult_result_T_74 ? 3'h4 : _GEN_763; // @[Jump.scala 155:19 186:26]
  wire  _GEN_797 = _execResult_result_T_74 ? 1'h0 : _GEN_761; // @[Jump.scala 155:19 152:20]
  wire [15:0] _GEN_798 = _execResult_result_T_74 ? operand : _GEN_762; // @[Jump.scala 155:19 153:20]
  wire  _GEN_800 = _execResult_result_T_74 ? 1'h0 : _GEN_777; // @[Jump.scala 146:17 155:19]
  wire [15:0] _GEN_801 = _execResult_result_T_22 ? execResult_result_result_19_memAddr : _GEN_778; // @[Jump.scala 155:19 170:24]
  wire [7:0] _GEN_802 = _execResult_result_T_22 ? regs_pc[7:0] : _GEN_779; // @[Jump.scala 155:19 171:24]
  wire [2:0] _GEN_817 = _execResult_result_T_22 ? 3'h3 : _GEN_796; // @[Jump.scala 155:19 175:26]
  wire  _GEN_820 = _execResult_result_T_22 ? 1'h0 : _GEN_797; // @[Jump.scala 155:19 152:20]
  wire [15:0] _GEN_821 = _execResult_result_T_22 ? operand : _GEN_798; // @[Jump.scala 155:19 153:20]
  wire  _GEN_823 = _execResult_result_T_22 ? 1'h0 : _GEN_800; // @[Jump.scala 146:17 155:19]
  wire [15:0] _GEN_824 = _execResult_result_T_21 ? execResult_result_result_19_memAddr : _GEN_801; // @[Jump.scala 155:19 162:24]
  wire [7:0] _GEN_825 = _execResult_result_T_21 ? regs_pc[15:8] : _GEN_802; // @[Jump.scala 155:19 163:24]
  wire  _GEN_826 = _execResult_result_T_21 | _GEN_633; // @[Jump.scala 155:19 164:25]
  wire [2:0] _GEN_840 = _execResult_result_T_21 ? 3'h2 : _GEN_817; // @[Jump.scala 155:19 167:26]
  wire  _GEN_843 = _execResult_result_T_21 ? 1'h0 : _GEN_820; // @[Jump.scala 155:19 152:20]
  wire [15:0] _GEN_844 = _execResult_result_T_21 ? operand : _GEN_821; // @[Jump.scala 155:19 153:20]
  wire  _GEN_846 = _execResult_result_T_21 ? 1'h0 : _GEN_823; // @[Jump.scala 146:17 155:19]
  wire [2:0] execResult_result_result_24_nextCycle = _execResult_result_T_20 ? 3'h1 : _GEN_840; // @[Jump.scala 155:19 159:26]
  wire [15:0] execResult_result_result_24_memAddr = _execResult_result_T_20 ? 16'h0 : _GEN_824; // @[Jump.scala 155:19 149:20]
  wire [7:0] execResult_result_result_24_memData = _execResult_result_T_20 ? 8'h0 : _GEN_825; // @[Jump.scala 155:19 150:20]
  wire  execResult_result_result_24_memWrite = _execResult_result_T_20 ? 1'h0 : _GEN_826; // @[Jump.scala 155:19 151:21]
  wire  execResult_result_result_24_memRead = _execResult_result_T_20 ? 1'h0 : _GEN_843; // @[Jump.scala 155:19 152:20]
  wire [15:0] execResult_result_result_24_operand = _execResult_result_T_20 ? operand : _GEN_844; // @[Jump.scala 155:19 153:20]
  wire  execResult_result_result_24_done = _execResult_result_T_20 ? 1'h0 : _GEN_846; // @[Jump.scala 146:17 155:19]
  wire [15:0] _GEN_872 = _execResult_result_T_74 ? _execResult_result_result_operand_T_4 : regs_pc; // @[Jump.scala 210:13 221:19 251:20]
  wire [7:0] _GEN_888 = _execResult_result_T_22 ? _execResult_result_newRegs_sp_T_3 : regs_sp; // @[Jump.scala 210:13 221:19 244:20]
  wire [7:0] _GEN_912 = _execResult_result_T_21 ? _execResult_result_newRegs_sp_T_3 : _GEN_888; // @[Jump.scala 221:19 236:20]
  wire [7:0] execResult_result_newRegs_24_sp = _execResult_result_T_20 ? _execResult_result_newRegs_sp_T_3 : _GEN_912; // @[Jump.scala 221:19 223:20]
  wire [15:0] _GEN_902 = _execResult_result_T_22 ? regs_pc : _GEN_872; // @[Jump.scala 210:13 221:19]
  wire [15:0] _GEN_927 = _execResult_result_T_21 ? regs_pc : _GEN_902; // @[Jump.scala 210:13 221:19]
  wire [15:0] execResult_result_newRegs_24_pc = _execResult_result_T_20 ? regs_pc : _GEN_927; // @[Jump.scala 210:13 221:19]
  wire  _GEN_906 = _execResult_result_T_21 ? io_memDataIn[0] : regs_flagC; // @[Jump.scala 210:13 221:19 230:23]
  wire  execResult_result_newRegs_24_flagC = _execResult_result_T_20 ? regs_flagC : _GEN_906; // @[Jump.scala 210:13 221:19]
  wire  _GEN_907 = _execResult_result_T_21 ? io_memDataIn[1] : regs_flagZ; // @[Jump.scala 210:13 221:19 231:23]
  wire  execResult_result_newRegs_24_flagZ = _execResult_result_T_20 ? regs_flagZ : _GEN_907; // @[Jump.scala 210:13 221:19]
  wire  _GEN_908 = _execResult_result_T_21 ? io_memDataIn[2] : regs_flagI; // @[Jump.scala 210:13 221:19 232:23]
  wire  execResult_result_newRegs_24_flagI = _execResult_result_T_20 ? regs_flagI : _GEN_908; // @[Jump.scala 210:13 221:19]
  wire  _GEN_909 = _execResult_result_T_21 ? io_memDataIn[3] : regs_flagD; // @[Jump.scala 210:13 221:19 233:23]
  wire  execResult_result_newRegs_24_flagD = _execResult_result_T_20 ? regs_flagD : _GEN_909; // @[Jump.scala 210:13 221:19]
  wire [15:0] _GEN_887 = _execResult_result_T_22 ? {{8'd0}, io_memDataIn} : operand; // @[Jump.scala 221:19 219:20 243:24]
  wire [15:0] _GEN_904 = _execResult_result_T_21 ? execResult_result_result_19_memAddr : _GEN_631; // @[Jump.scala 221:19 228:24]
  wire [15:0] _GEN_926 = _execResult_result_T_21 ? operand : _GEN_887; // @[Jump.scala 221:19 219:20]
  wire [15:0] execResult_result_result_25_memAddr = _execResult_result_T_20 ? 16'h0 : _GEN_904; // @[Jump.scala 221:19 215:20]
  wire [15:0] execResult_result_result_25_operand = _execResult_result_T_20 ? operand : _GEN_926; // @[Jump.scala 221:19 219:20]
  wire  _GEN_954 = 8'h40 == opcode & execResult_result_result_22_done; // @[CPU6502Core.scala 89:20 189:27 87:12]
  wire [2:0] _GEN_955 = 8'h40 == opcode ? execResult_result_result_22_nextCycle : 3'h0; // @[CPU6502Core.scala 89:20 189:27 87:12]
  wire [7:0] _GEN_959 = 8'h40 == opcode ? execResult_result_newRegs_24_sp : regs_sp; // @[CPU6502Core.scala 89:20 189:27 87:12]
  wire [15:0] _GEN_960 = 8'h40 == opcode ? execResult_result_newRegs_24_pc : regs_pc; // @[CPU6502Core.scala 89:20 189:27 87:12]
  wire  _GEN_961 = 8'h40 == opcode ? execResult_result_newRegs_24_flagC : regs_flagC; // @[CPU6502Core.scala 89:20 189:27 87:12]
  wire  _GEN_962 = 8'h40 == opcode ? execResult_result_newRegs_24_flagZ : regs_flagZ; // @[CPU6502Core.scala 89:20 189:27 87:12]
  wire  _GEN_963 = 8'h40 == opcode ? execResult_result_newRegs_24_flagI : regs_flagI; // @[CPU6502Core.scala 89:20 189:27 87:12]
  wire  _GEN_964 = 8'h40 == opcode ? execResult_result_newRegs_24_flagD : regs_flagD; // @[CPU6502Core.scala 89:20 189:27 87:12]
  wire  _GEN_966 = 8'h40 == opcode ? execResult_result_newRegs_7_flagV : regs_flagV; // @[CPU6502Core.scala 89:20 189:27 87:12]
  wire  _GEN_967 = 8'h40 == opcode ? execResult_result_newRegs_7_flagN : regs_flagN; // @[CPU6502Core.scala 89:20 189:27 87:12]
  wire [15:0] _GEN_968 = 8'h40 == opcode ? execResult_result_result_25_memAddr : 16'h0; // @[CPU6502Core.scala 89:20 189:27 87:12]
  wire  _GEN_971 = 8'h40 == opcode & execResult_result_result_24_memWrite; // @[CPU6502Core.scala 89:20 189:27 87:12]
  wire [15:0] _GEN_972 = 8'h40 == opcode ? execResult_result_result_25_operand : operand; // @[CPU6502Core.scala 89:20 189:27 87:12]
  wire  _GEN_973 = 8'h0 == opcode ? execResult_result_result_24_done : _GEN_954; // @[CPU6502Core.scala 89:20 188:27]
  wire [2:0] _GEN_974 = 8'h0 == opcode ? execResult_result_result_24_nextCycle : _GEN_955; // @[CPU6502Core.scala 89:20 188:27]
  wire [7:0] _GEN_978 = 8'h0 == opcode ? execResult_result_newRegs_23_sp : _GEN_959; // @[CPU6502Core.scala 89:20 188:27]
  wire [15:0] _GEN_979 = 8'h0 == opcode ? execResult_result_newRegs_23_pc : _GEN_960; // @[CPU6502Core.scala 89:20 188:27]
  wire  _GEN_980 = 8'h0 == opcode ? regs_flagC : _GEN_961; // @[CPU6502Core.scala 89:20 188:27]
  wire  _GEN_981 = 8'h0 == opcode ? regs_flagZ : _GEN_962; // @[CPU6502Core.scala 89:20 188:27]
  wire  _GEN_982 = 8'h0 == opcode ? execResult_result_newRegs_23_flagI : _GEN_963; // @[CPU6502Core.scala 89:20 188:27]
  wire  _GEN_983 = 8'h0 == opcode ? regs_flagD : _GEN_964; // @[CPU6502Core.scala 89:20 188:27]
  wire  _GEN_985 = 8'h0 == opcode ? regs_flagV : _GEN_966; // @[CPU6502Core.scala 89:20 188:27]
  wire  _GEN_986 = 8'h0 == opcode ? regs_flagN : _GEN_967; // @[CPU6502Core.scala 89:20 188:27]
  wire [15:0] _GEN_987 = 8'h0 == opcode ? execResult_result_result_24_memAddr : _GEN_968; // @[CPU6502Core.scala 89:20 188:27]
  wire [7:0] _GEN_988 = 8'h0 == opcode ? execResult_result_result_24_memData : 8'h0; // @[CPU6502Core.scala 89:20 188:27]
  wire  _GEN_989 = 8'h0 == opcode & execResult_result_result_24_memWrite; // @[CPU6502Core.scala 89:20 188:27]
  wire  _GEN_990 = 8'h0 == opcode ? execResult_result_result_24_memRead : _GEN_971; // @[CPU6502Core.scala 89:20 188:27]
  wire [15:0] _GEN_991 = 8'h0 == opcode ? execResult_result_result_24_operand : _GEN_972; // @[CPU6502Core.scala 89:20 188:27]
  wire  _GEN_992 = 8'h60 == opcode ? execResult_result_result_6_done : _GEN_973; // @[CPU6502Core.scala 89:20 187:27]
  wire [2:0] _GEN_993 = 8'h60 == opcode ? execResult_result_result_6_nextCycle : _GEN_974; // @[CPU6502Core.scala 89:20 187:27]
  wire [7:0] _GEN_997 = 8'h60 == opcode ? execResult_result_newRegs_22_sp : _GEN_978; // @[CPU6502Core.scala 89:20 187:27]
  wire [15:0] _GEN_998 = 8'h60 == opcode ? execResult_result_newRegs_22_pc : _GEN_979; // @[CPU6502Core.scala 89:20 187:27]
  wire  _GEN_999 = 8'h60 == opcode ? regs_flagC : _GEN_980; // @[CPU6502Core.scala 89:20 187:27]
  wire  _GEN_1000 = 8'h60 == opcode ? regs_flagZ : _GEN_981; // @[CPU6502Core.scala 89:20 187:27]
  wire  _GEN_1001 = 8'h60 == opcode ? regs_flagI : _GEN_982; // @[CPU6502Core.scala 89:20 187:27]
  wire  _GEN_1002 = 8'h60 == opcode ? regs_flagD : _GEN_983; // @[CPU6502Core.scala 89:20 187:27]
  wire  _GEN_1004 = 8'h60 == opcode ? regs_flagV : _GEN_985; // @[CPU6502Core.scala 89:20 187:27]
  wire  _GEN_1005 = 8'h60 == opcode ? regs_flagN : _GEN_986; // @[CPU6502Core.scala 89:20 187:27]
  wire [15:0] _GEN_1006 = 8'h60 == opcode ? execResult_result_result_23_memAddr : _GEN_987; // @[CPU6502Core.scala 89:20 187:27]
  wire [7:0] _GEN_1007 = 8'h60 == opcode ? 8'h0 : _GEN_988; // @[CPU6502Core.scala 89:20 187:27]
  wire  _GEN_1008 = 8'h60 == opcode ? 1'h0 : _GEN_989; // @[CPU6502Core.scala 89:20 187:27]
  wire  _GEN_1009 = 8'h60 == opcode ? execResult_result_result_23_memRead : _GEN_990; // @[CPU6502Core.scala 89:20 187:27]
  wire [15:0] _GEN_1010 = 8'h60 == opcode ? execResult_result_result_23_operand : _GEN_991; // @[CPU6502Core.scala 89:20 187:27]
  wire  _GEN_1011 = 8'h20 == opcode ? execResult_result_result_22_done : _GEN_992; // @[CPU6502Core.scala 89:20 186:27]
  wire [2:0] _GEN_1012 = 8'h20 == opcode ? execResult_result_result_22_nextCycle : _GEN_993; // @[CPU6502Core.scala 89:20 186:27]
  wire [7:0] _GEN_1016 = 8'h20 == opcode ? execResult_result_newRegs_21_sp : _GEN_997; // @[CPU6502Core.scala 89:20 186:27]
  wire [15:0] _GEN_1017 = 8'h20 == opcode ? execResult_result_newRegs_21_pc : _GEN_998; // @[CPU6502Core.scala 89:20 186:27]
  wire  _GEN_1018 = 8'h20 == opcode ? regs_flagC : _GEN_999; // @[CPU6502Core.scala 89:20 186:27]
  wire  _GEN_1019 = 8'h20 == opcode ? regs_flagZ : _GEN_1000; // @[CPU6502Core.scala 89:20 186:27]
  wire  _GEN_1020 = 8'h20 == opcode ? regs_flagI : _GEN_1001; // @[CPU6502Core.scala 89:20 186:27]
  wire  _GEN_1021 = 8'h20 == opcode ? regs_flagD : _GEN_1002; // @[CPU6502Core.scala 89:20 186:27]
  wire  _GEN_1023 = 8'h20 == opcode ? regs_flagV : _GEN_1004; // @[CPU6502Core.scala 89:20 186:27]
  wire  _GEN_1024 = 8'h20 == opcode ? regs_flagN : _GEN_1005; // @[CPU6502Core.scala 89:20 186:27]
  wire [15:0] _GEN_1025 = 8'h20 == opcode ? execResult_result_result_22_memAddr : _GEN_1006; // @[CPU6502Core.scala 89:20 186:27]
  wire [7:0] _GEN_1026 = 8'h20 == opcode ? execResult_result_result_22_memData : _GEN_1007; // @[CPU6502Core.scala 89:20 186:27]
  wire  _GEN_1027 = 8'h20 == opcode ? execResult_result_result_22_memWrite : _GEN_1008; // @[CPU6502Core.scala 89:20 186:27]
  wire  _GEN_1028 = 8'h20 == opcode ? execResult_result_result_6_memRead : _GEN_1009; // @[CPU6502Core.scala 89:20 186:27]
  wire [15:0] _GEN_1029 = 8'h20 == opcode ? execResult_result_result_17_operand : _GEN_1010; // @[CPU6502Core.scala 89:20 186:27]
  wire  _GEN_1030 = 8'h4c == opcode ? execResult_result_result_8_done : _GEN_1011; // @[CPU6502Core.scala 89:20 185:27]
  wire [2:0] _GEN_1031 = 8'h4c == opcode ? execResult_result_result_8_nextCycle : _GEN_1012; // @[CPU6502Core.scala 89:20 185:27]
  wire [7:0] _GEN_1035 = 8'h4c == opcode ? regs_sp : _GEN_1016; // @[CPU6502Core.scala 89:20 185:27]
  wire [15:0] _GEN_1036 = 8'h4c == opcode ? execResult_result_newRegs_20_pc : _GEN_1017; // @[CPU6502Core.scala 89:20 185:27]
  wire  _GEN_1037 = 8'h4c == opcode ? regs_flagC : _GEN_1018; // @[CPU6502Core.scala 89:20 185:27]
  wire  _GEN_1038 = 8'h4c == opcode ? regs_flagZ : _GEN_1019; // @[CPU6502Core.scala 89:20 185:27]
  wire  _GEN_1039 = 8'h4c == opcode ? regs_flagI : _GEN_1020; // @[CPU6502Core.scala 89:20 185:27]
  wire  _GEN_1040 = 8'h4c == opcode ? regs_flagD : _GEN_1021; // @[CPU6502Core.scala 89:20 185:27]
  wire  _GEN_1042 = 8'h4c == opcode ? regs_flagV : _GEN_1023; // @[CPU6502Core.scala 89:20 185:27]
  wire  _GEN_1043 = 8'h4c == opcode ? regs_flagN : _GEN_1024; // @[CPU6502Core.scala 89:20 185:27]
  wire [15:0] _GEN_1044 = 8'h4c == opcode ? execResult_result_result_21_memAddr : _GEN_1025; // @[CPU6502Core.scala 89:20 185:27]
  wire [7:0] _GEN_1045 = 8'h4c == opcode ? 8'h0 : _GEN_1026; // @[CPU6502Core.scala 89:20 185:27]
  wire  _GEN_1046 = 8'h4c == opcode ? 1'h0 : _GEN_1027; // @[CPU6502Core.scala 89:20 185:27]
  wire  _GEN_1047 = 8'h4c == opcode ? execResult_result_result_6_memRead : _GEN_1028; // @[CPU6502Core.scala 89:20 185:27]
  wire [15:0] _GEN_1048 = 8'h4c == opcode ? execResult_result_result_6_operand : _GEN_1029; // @[CPU6502Core.scala 89:20 185:27]
  wire  _GEN_1049 = 8'h68 == opcode | 8'h28 == opcode ? execResult_result_result_8_done : _GEN_1030; // @[CPU6502Core.scala 181:16 89:20]
  wire [2:0] _GEN_1050 = 8'h68 == opcode | 8'h28 == opcode ? execResult_result_result_8_nextCycle : _GEN_1031; // @[CPU6502Core.scala 181:16 89:20]
  wire [7:0] _GEN_1051 = 8'h68 == opcode | 8'h28 == opcode ? execResult_result_newRegs_19_a : regs_a; // @[CPU6502Core.scala 181:16 89:20]
  wire [7:0] _GEN_1054 = 8'h68 == opcode | 8'h28 == opcode ? execResult_result_newRegs_19_sp : _GEN_1035; // @[CPU6502Core.scala 181:16 89:20]
  wire [15:0] _GEN_1055 = 8'h68 == opcode | 8'h28 == opcode ? regs_pc : _GEN_1036; // @[CPU6502Core.scala 181:16 89:20]
  wire  _GEN_1056 = 8'h68 == opcode | 8'h28 == opcode ? execResult_result_newRegs_19_flagC : _GEN_1037; // @[CPU6502Core.scala 181:16 89:20]
  wire  _GEN_1057 = 8'h68 == opcode | 8'h28 == opcode ? execResult_result_newRegs_19_flagZ : _GEN_1038; // @[CPU6502Core.scala 181:16 89:20]
  wire  _GEN_1058 = 8'h68 == opcode | 8'h28 == opcode ? execResult_result_newRegs_19_flagI : _GEN_1039; // @[CPU6502Core.scala 181:16 89:20]
  wire  _GEN_1059 = 8'h68 == opcode | 8'h28 == opcode ? execResult_result_newRegs_19_flagD : _GEN_1040; // @[CPU6502Core.scala 181:16 89:20]
  wire  _GEN_1061 = 8'h68 == opcode | 8'h28 == opcode ? execResult_result_newRegs_19_flagV : _GEN_1042; // @[CPU6502Core.scala 181:16 89:20]
  wire  _GEN_1062 = 8'h68 == opcode | 8'h28 == opcode ? execResult_result_newRegs_19_flagN : _GEN_1043; // @[CPU6502Core.scala 181:16 89:20]
  wire [15:0] _GEN_1063 = 8'h68 == opcode | 8'h28 == opcode ? execResult_result_result_20_memAddr : _GEN_1044; // @[CPU6502Core.scala 181:16 89:20]
  wire [7:0] _GEN_1064 = 8'h68 == opcode | 8'h28 == opcode ? 8'h0 : _GEN_1045; // @[CPU6502Core.scala 181:16 89:20]
  wire  _GEN_1065 = 8'h68 == opcode | 8'h28 == opcode ? 1'h0 : _GEN_1046; // @[CPU6502Core.scala 181:16 89:20]
  wire  _GEN_1066 = 8'h68 == opcode | 8'h28 == opcode ? execResult_result_result_8_done : _GEN_1047; // @[CPU6502Core.scala 181:16 89:20]
  wire [15:0] _GEN_1067 = 8'h68 == opcode | 8'h28 == opcode ? 16'h0 : _GEN_1048; // @[CPU6502Core.scala 181:16 89:20]
  wire  _GEN_1068 = 8'h48 == opcode | 8'h8 == opcode | _GEN_1049; // @[CPU6502Core.scala 176:16 89:20]
  wire [2:0] _GEN_1069 = 8'h48 == opcode | 8'h8 == opcode ? 3'h0 : _GEN_1050; // @[CPU6502Core.scala 176:16 89:20]
  wire [7:0] _GEN_1070 = 8'h48 == opcode | 8'h8 == opcode ? regs_a : _GEN_1051; // @[CPU6502Core.scala 176:16 89:20]
  wire [7:0] _GEN_1073 = 8'h48 == opcode | 8'h8 == opcode ? execResult_result_newRegs_18_sp : _GEN_1054; // @[CPU6502Core.scala 176:16 89:20]
  wire [15:0] _GEN_1074 = 8'h48 == opcode | 8'h8 == opcode ? regs_pc : _GEN_1055; // @[CPU6502Core.scala 176:16 89:20]
  wire  _GEN_1075 = 8'h48 == opcode | 8'h8 == opcode ? regs_flagC : _GEN_1056; // @[CPU6502Core.scala 176:16 89:20]
  wire  _GEN_1076 = 8'h48 == opcode | 8'h8 == opcode ? regs_flagZ : _GEN_1057; // @[CPU6502Core.scala 176:16 89:20]
  wire  _GEN_1077 = 8'h48 == opcode | 8'h8 == opcode ? regs_flagI : _GEN_1058; // @[CPU6502Core.scala 176:16 89:20]
  wire  _GEN_1078 = 8'h48 == opcode | 8'h8 == opcode ? regs_flagD : _GEN_1059; // @[CPU6502Core.scala 176:16 89:20]
  wire  _GEN_1080 = 8'h48 == opcode | 8'h8 == opcode ? regs_flagV : _GEN_1061; // @[CPU6502Core.scala 176:16 89:20]
  wire  _GEN_1081 = 8'h48 == opcode | 8'h8 == opcode ? regs_flagN : _GEN_1062; // @[CPU6502Core.scala 176:16 89:20]
  wire [15:0] _GEN_1082 = 8'h48 == opcode | 8'h8 == opcode ? execResult_result_result_19_memAddr : _GEN_1063; // @[CPU6502Core.scala 176:16 89:20]
  wire [7:0] _GEN_1083 = 8'h48 == opcode | 8'h8 == opcode ? execResult_result_pushData : _GEN_1064; // @[CPU6502Core.scala 176:16 89:20]
  wire  _GEN_1084 = 8'h48 == opcode | 8'h8 == opcode | _GEN_1065; // @[CPU6502Core.scala 176:16 89:20]
  wire  _GEN_1085 = 8'h48 == opcode | 8'h8 == opcode ? 1'h0 : _GEN_1066; // @[CPU6502Core.scala 176:16 89:20]
  wire [15:0] _GEN_1086 = 8'h48 == opcode | 8'h8 == opcode ? 16'h0 : _GEN_1067; // @[CPU6502Core.scala 176:16 89:20]
  wire  _GEN_1087 = 8'hbd == opcode | 8'hb9 == opcode ? execResult_result_result_6_done : _GEN_1068; // @[CPU6502Core.scala 171:16 89:20]
  wire [2:0] _GEN_1088 = 8'hbd == opcode | 8'hb9 == opcode ? execResult_result_result_6_nextCycle : _GEN_1069; // @[CPU6502Core.scala 171:16 89:20]
  wire [7:0] _GEN_1089 = 8'hbd == opcode | 8'hb9 == opcode ? execResult_result_newRegs_17_a : _GEN_1070; // @[CPU6502Core.scala 171:16 89:20]
  wire [7:0] _GEN_1092 = 8'hbd == opcode | 8'hb9 == opcode ? regs_sp : _GEN_1073; // @[CPU6502Core.scala 171:16 89:20]
  wire [15:0] _GEN_1093 = 8'hbd == opcode | 8'hb9 == opcode ? execResult_result_newRegs_16_pc : _GEN_1074; // @[CPU6502Core.scala 171:16 89:20]
  wire  _GEN_1094 = 8'hbd == opcode | 8'hb9 == opcode ? regs_flagC : _GEN_1075; // @[CPU6502Core.scala 171:16 89:20]
  wire  _GEN_1095 = 8'hbd == opcode | 8'hb9 == opcode ? execResult_result_newRegs_17_flagZ : _GEN_1076; // @[CPU6502Core.scala 171:16 89:20]
  wire  _GEN_1096 = 8'hbd == opcode | 8'hb9 == opcode ? regs_flagI : _GEN_1077; // @[CPU6502Core.scala 171:16 89:20]
  wire  _GEN_1097 = 8'hbd == opcode | 8'hb9 == opcode ? regs_flagD : _GEN_1078; // @[CPU6502Core.scala 171:16 89:20]
  wire  _GEN_1099 = 8'hbd == opcode | 8'hb9 == opcode ? regs_flagV : _GEN_1080; // @[CPU6502Core.scala 171:16 89:20]
  wire  _GEN_1100 = 8'hbd == opcode | 8'hb9 == opcode ? execResult_result_newRegs_17_flagN : _GEN_1081; // @[CPU6502Core.scala 171:16 89:20]
  wire [15:0] _GEN_1101 = 8'hbd == opcode | 8'hb9 == opcode ? execResult_result_result_17_memAddr : _GEN_1082; // @[CPU6502Core.scala 171:16 89:20]
  wire [7:0] _GEN_1102 = 8'hbd == opcode | 8'hb9 == opcode ? 8'h0 : _GEN_1083; // @[CPU6502Core.scala 171:16 89:20]
  wire  _GEN_1103 = 8'hbd == opcode | 8'hb9 == opcode ? 1'h0 : _GEN_1084; // @[CPU6502Core.scala 171:16 89:20]
  wire  _GEN_1104 = 8'hbd == opcode | 8'hb9 == opcode ? execResult_result_result_18_memRead : _GEN_1085; // @[CPU6502Core.scala 171:16 89:20]
  wire [15:0] _GEN_1105 = 8'hbd == opcode | 8'hb9 == opcode ? execResult_result_result_18_operand : _GEN_1086; // @[CPU6502Core.scala 171:16 89:20]
  wire  _GEN_1106 = 8'had == opcode | 8'h8d == opcode ? execResult_result_result_6_done : _GEN_1087; // @[CPU6502Core.scala 166:16 89:20]
  wire [2:0] _GEN_1107 = 8'had == opcode | 8'h8d == opcode ? execResult_result_result_6_nextCycle : _GEN_1088; // @[CPU6502Core.scala 166:16 89:20]
  wire [7:0] _GEN_1108 = 8'had == opcode | 8'h8d == opcode ? execResult_result_newRegs_16_a : _GEN_1089; // @[CPU6502Core.scala 166:16 89:20]
  wire [7:0] _GEN_1111 = 8'had == opcode | 8'h8d == opcode ? regs_sp : _GEN_1092; // @[CPU6502Core.scala 166:16 89:20]
  wire [15:0] _GEN_1112 = 8'had == opcode | 8'h8d == opcode ? execResult_result_newRegs_16_pc : _GEN_1093; // @[CPU6502Core.scala 166:16 89:20]
  wire  _GEN_1113 = 8'had == opcode | 8'h8d == opcode ? regs_flagC : _GEN_1094; // @[CPU6502Core.scala 166:16 89:20]
  wire  _GEN_1114 = 8'had == opcode | 8'h8d == opcode ? execResult_result_newRegs_16_flagZ : _GEN_1095; // @[CPU6502Core.scala 166:16 89:20]
  wire  _GEN_1115 = 8'had == opcode | 8'h8d == opcode ? regs_flagI : _GEN_1096; // @[CPU6502Core.scala 166:16 89:20]
  wire  _GEN_1116 = 8'had == opcode | 8'h8d == opcode ? regs_flagD : _GEN_1097; // @[CPU6502Core.scala 166:16 89:20]
  wire  _GEN_1118 = 8'had == opcode | 8'h8d == opcode ? regs_flagV : _GEN_1099; // @[CPU6502Core.scala 166:16 89:20]
  wire  _GEN_1119 = 8'had == opcode | 8'h8d == opcode ? execResult_result_newRegs_16_flagN : _GEN_1100; // @[CPU6502Core.scala 166:16 89:20]
  wire [15:0] _GEN_1120 = 8'had == opcode | 8'h8d == opcode ? execResult_result_result_17_memAddr : _GEN_1101; // @[CPU6502Core.scala 166:16 89:20]
  wire [7:0] _GEN_1121 = 8'had == opcode | 8'h8d == opcode ? execResult_result_result_17_memData : _GEN_1102; // @[CPU6502Core.scala 166:16 89:20]
  wire  _GEN_1122 = 8'had == opcode | 8'h8d == opcode ? execResult_result_result_17_memWrite : _GEN_1103; // @[CPU6502Core.scala 166:16 89:20]
  wire  _GEN_1123 = 8'had == opcode | 8'h8d == opcode ? execResult_result_result_17_memRead : _GEN_1104; // @[CPU6502Core.scala 166:16 89:20]
  wire [15:0] _GEN_1124 = 8'had == opcode | 8'h8d == opcode ? execResult_result_result_17_operand : _GEN_1105; // @[CPU6502Core.scala 166:16 89:20]
  wire  _GEN_1125 = 8'hb5 == opcode | 8'h95 == opcode ? execResult_result_result_8_done : _GEN_1106; // @[CPU6502Core.scala 161:16 89:20]
  wire [2:0] _GEN_1126 = 8'hb5 == opcode | 8'h95 == opcode ? execResult_result_result_8_nextCycle : _GEN_1107; // @[CPU6502Core.scala 161:16 89:20]
  wire [7:0] _GEN_1127 = 8'hb5 == opcode | 8'h95 == opcode ? execResult_result_newRegs_15_a : _GEN_1108; // @[CPU6502Core.scala 161:16 89:20]
  wire [7:0] _GEN_1130 = 8'hb5 == opcode | 8'h95 == opcode ? regs_sp : _GEN_1111; // @[CPU6502Core.scala 161:16 89:20]
  wire [15:0] _GEN_1131 = 8'hb5 == opcode | 8'h95 == opcode ? execResult_result_newRegs_5_pc : _GEN_1112; // @[CPU6502Core.scala 161:16 89:20]
  wire  _GEN_1132 = 8'hb5 == opcode | 8'h95 == opcode ? regs_flagC : _GEN_1113; // @[CPU6502Core.scala 161:16 89:20]
  wire  _GEN_1133 = 8'hb5 == opcode | 8'h95 == opcode ? execResult_result_newRegs_15_flagZ : _GEN_1114; // @[CPU6502Core.scala 161:16 89:20]
  wire  _GEN_1134 = 8'hb5 == opcode | 8'h95 == opcode ? regs_flagI : _GEN_1115; // @[CPU6502Core.scala 161:16 89:20]
  wire  _GEN_1135 = 8'hb5 == opcode | 8'h95 == opcode ? regs_flagD : _GEN_1116; // @[CPU6502Core.scala 161:16 89:20]
  wire  _GEN_1137 = 8'hb5 == opcode | 8'h95 == opcode ? regs_flagV : _GEN_1118; // @[CPU6502Core.scala 161:16 89:20]
  wire  _GEN_1138 = 8'hb5 == opcode | 8'h95 == opcode ? execResult_result_newRegs_15_flagN : _GEN_1119; // @[CPU6502Core.scala 161:16 89:20]
  wire [15:0] _GEN_1139 = 8'hb5 == opcode | 8'h95 == opcode ? execResult_result_result_8_memAddr : _GEN_1120; // @[CPU6502Core.scala 161:16 89:20]
  wire [7:0] _GEN_1140 = 8'hb5 == opcode | 8'h95 == opcode ? execResult_result_result_16_memData : _GEN_1121; // @[CPU6502Core.scala 161:16 89:20]
  wire  _GEN_1141 = 8'hb5 == opcode | 8'h95 == opcode ? execResult_result_result_16_memWrite : _GEN_1122; // @[CPU6502Core.scala 161:16 89:20]
  wire  _GEN_1142 = 8'hb5 == opcode | 8'h95 == opcode ? execResult_result_result_16_memRead : _GEN_1123; // @[CPU6502Core.scala 161:16 89:20]
  wire [15:0] _GEN_1143 = 8'hb5 == opcode | 8'h95 == opcode ? execResult_result_result_16_operand : _GEN_1124; // @[CPU6502Core.scala 161:16 89:20]
  wire  _GEN_1144 = 8'ha5 == opcode | 8'h85 == opcode | 8'h86 == opcode | 8'h84 == opcode ?
    execResult_result_result_8_done : _GEN_1125; // @[CPU6502Core.scala 156:16 89:20]
  wire [2:0] _GEN_1145 = 8'ha5 == opcode | 8'h85 == opcode | 8'h86 == opcode | 8'h84 == opcode ?
    execResult_result_result_8_nextCycle : _GEN_1126; // @[CPU6502Core.scala 156:16 89:20]
  wire [7:0] _GEN_1146 = 8'ha5 == opcode | 8'h85 == opcode | 8'h86 == opcode | 8'h84 == opcode ?
    execResult_result_newRegs_14_a : _GEN_1127; // @[CPU6502Core.scala 156:16 89:20]
  wire [7:0] _GEN_1149 = 8'ha5 == opcode | 8'h85 == opcode | 8'h86 == opcode | 8'h84 == opcode ? regs_sp : _GEN_1130; // @[CPU6502Core.scala 156:16 89:20]
  wire [15:0] _GEN_1150 = 8'ha5 == opcode | 8'h85 == opcode | 8'h86 == opcode | 8'h84 == opcode ?
    execResult_result_newRegs_5_pc : _GEN_1131; // @[CPU6502Core.scala 156:16 89:20]
  wire  _GEN_1151 = 8'ha5 == opcode | 8'h85 == opcode | 8'h86 == opcode | 8'h84 == opcode ? regs_flagC : _GEN_1132; // @[CPU6502Core.scala 156:16 89:20]
  wire  _GEN_1152 = 8'ha5 == opcode | 8'h85 == opcode | 8'h86 == opcode | 8'h84 == opcode ?
    execResult_result_newRegs_14_flagZ : _GEN_1133; // @[CPU6502Core.scala 156:16 89:20]
  wire  _GEN_1153 = 8'ha5 == opcode | 8'h85 == opcode | 8'h86 == opcode | 8'h84 == opcode ? regs_flagI : _GEN_1134; // @[CPU6502Core.scala 156:16 89:20]
  wire  _GEN_1154 = 8'ha5 == opcode | 8'h85 == opcode | 8'h86 == opcode | 8'h84 == opcode ? regs_flagD : _GEN_1135; // @[CPU6502Core.scala 156:16 89:20]
  wire  _GEN_1156 = 8'ha5 == opcode | 8'h85 == opcode | 8'h86 == opcode | 8'h84 == opcode ? regs_flagV : _GEN_1137; // @[CPU6502Core.scala 156:16 89:20]
  wire  _GEN_1157 = 8'ha5 == opcode | 8'h85 == opcode | 8'h86 == opcode | 8'h84 == opcode ?
    execResult_result_newRegs_14_flagN : _GEN_1138; // @[CPU6502Core.scala 156:16 89:20]
  wire [15:0] _GEN_1158 = 8'ha5 == opcode | 8'h85 == opcode | 8'h86 == opcode | 8'h84 == opcode ?
    execResult_result_result_8_memAddr : _GEN_1139; // @[CPU6502Core.scala 156:16 89:20]
  wire [7:0] _GEN_1159 = 8'ha5 == opcode | 8'h85 == opcode | 8'h86 == opcode | 8'h84 == opcode ?
    execResult_result_result_15_memData : _GEN_1140; // @[CPU6502Core.scala 156:16 89:20]
  wire  _GEN_1160 = 8'ha5 == opcode | 8'h85 == opcode | 8'h86 == opcode | 8'h84 == opcode ?
    execResult_result_result_15_memWrite : _GEN_1141; // @[CPU6502Core.scala 156:16 89:20]
  wire  _GEN_1161 = 8'ha5 == opcode | 8'h85 == opcode | 8'h86 == opcode | 8'h84 == opcode ?
    execResult_result_result_15_memRead : _GEN_1142; // @[CPU6502Core.scala 156:16 89:20]
  wire [15:0] _GEN_1162 = 8'ha5 == opcode | 8'h85 == opcode | 8'h86 == opcode | 8'h84 == opcode ?
    execResult_result_result_6_operand : _GEN_1143; // @[CPU6502Core.scala 156:16 89:20]
  wire  _GEN_1163 = 8'ha9 == opcode | 8'ha2 == opcode | 8'ha0 == opcode | _GEN_1144; // @[CPU6502Core.scala 151:16 89:20]
  wire [2:0] _GEN_1164 = 8'ha9 == opcode | 8'ha2 == opcode | 8'ha0 == opcode ? 3'h0 : _GEN_1145; // @[CPU6502Core.scala 151:16 89:20]
  wire [7:0] _GEN_1165 = 8'ha9 == opcode | 8'ha2 == opcode | 8'ha0 == opcode ? execResult_result_newRegs_13_a :
    _GEN_1146; // @[CPU6502Core.scala 151:16 89:20]
  wire [7:0] _GEN_1166 = 8'ha9 == opcode | 8'ha2 == opcode | 8'ha0 == opcode ? execResult_result_newRegs_13_x : regs_x; // @[CPU6502Core.scala 151:16 89:20]
  wire [7:0] _GEN_1167 = 8'ha9 == opcode | 8'ha2 == opcode | 8'ha0 == opcode ? execResult_result_newRegs_13_y : regs_y; // @[CPU6502Core.scala 151:16 89:20]
  wire [7:0] _GEN_1168 = 8'ha9 == opcode | 8'ha2 == opcode | 8'ha0 == opcode ? regs_sp : _GEN_1149; // @[CPU6502Core.scala 151:16 89:20]
  wire [15:0] _GEN_1169 = 8'ha9 == opcode | 8'ha2 == opcode | 8'ha0 == opcode ? _regs_pc_T_1 : _GEN_1150; // @[CPU6502Core.scala 151:16 89:20]
  wire  _GEN_1170 = 8'ha9 == opcode | 8'ha2 == opcode | 8'ha0 == opcode ? regs_flagC : _GEN_1151; // @[CPU6502Core.scala 151:16 89:20]
  wire  _GEN_1171 = 8'ha9 == opcode | 8'ha2 == opcode | 8'ha0 == opcode ? execResult_result_newRegs_13_flagZ : _GEN_1152
    ; // @[CPU6502Core.scala 151:16 89:20]
  wire  _GEN_1172 = 8'ha9 == opcode | 8'ha2 == opcode | 8'ha0 == opcode ? regs_flagI : _GEN_1153; // @[CPU6502Core.scala 151:16 89:20]
  wire  _GEN_1173 = 8'ha9 == opcode | 8'ha2 == opcode | 8'ha0 == opcode ? regs_flagD : _GEN_1154; // @[CPU6502Core.scala 151:16 89:20]
  wire  _GEN_1175 = 8'ha9 == opcode | 8'ha2 == opcode | 8'ha0 == opcode ? regs_flagV : _GEN_1156; // @[CPU6502Core.scala 151:16 89:20]
  wire  _GEN_1176 = 8'ha9 == opcode | 8'ha2 == opcode | 8'ha0 == opcode ? io_memDataIn[7] : _GEN_1157; // @[CPU6502Core.scala 151:16 89:20]
  wire [15:0] _GEN_1177 = 8'ha9 == opcode | 8'ha2 == opcode | 8'ha0 == opcode ? regs_pc : _GEN_1158; // @[CPU6502Core.scala 151:16 89:20]
  wire [7:0] _GEN_1178 = 8'ha9 == opcode | 8'ha2 == opcode | 8'ha0 == opcode ? 8'h0 : _GEN_1159; // @[CPU6502Core.scala 151:16 89:20]
  wire  _GEN_1179 = 8'ha9 == opcode | 8'ha2 == opcode | 8'ha0 == opcode ? 1'h0 : _GEN_1160; // @[CPU6502Core.scala 151:16 89:20]
  wire  _GEN_1180 = 8'ha9 == opcode | 8'ha2 == opcode | 8'ha0 == opcode | _GEN_1161; // @[CPU6502Core.scala 151:16 89:20]
  wire [15:0] _GEN_1181 = 8'ha9 == opcode | 8'ha2 == opcode | 8'ha0 == opcode ? 16'h0 : _GEN_1162; // @[CPU6502Core.scala 151:16 89:20]
  wire  _GEN_1182 = 8'hf0 == opcode | 8'hd0 == opcode | 8'hb0 == opcode | 8'h90 == opcode | 8'h30 == opcode | 8'h10 ==
    opcode | 8'h50 == opcode | 8'h70 == opcode | _GEN_1163; // @[CPU6502Core.scala 146:16 89:20]
  wire [2:0] _GEN_1183 = 8'hf0 == opcode | 8'hd0 == opcode | 8'hb0 == opcode | 8'h90 == opcode | 8'h30 == opcode | 8'h10
     == opcode | 8'h50 == opcode | 8'h70 == opcode ? 3'h0 : _GEN_1164; // @[CPU6502Core.scala 146:16 89:20]
  wire [7:0] _GEN_1184 = 8'hf0 == opcode | 8'hd0 == opcode | 8'hb0 == opcode | 8'h90 == opcode | 8'h30 == opcode | 8'h10
     == opcode | 8'h50 == opcode | 8'h70 == opcode ? regs_a : _GEN_1165; // @[CPU6502Core.scala 146:16 89:20]
  wire [7:0] _GEN_1185 = 8'hf0 == opcode | 8'hd0 == opcode | 8'hb0 == opcode | 8'h90 == opcode | 8'h30 == opcode | 8'h10
     == opcode | 8'h50 == opcode | 8'h70 == opcode ? regs_x : _GEN_1166; // @[CPU6502Core.scala 146:16 89:20]
  wire [7:0] _GEN_1186 = 8'hf0 == opcode | 8'hd0 == opcode | 8'hb0 == opcode | 8'h90 == opcode | 8'h30 == opcode | 8'h10
     == opcode | 8'h50 == opcode | 8'h70 == opcode ? regs_y : _GEN_1167; // @[CPU6502Core.scala 146:16 89:20]
  wire [7:0] _GEN_1187 = 8'hf0 == opcode | 8'hd0 == opcode | 8'hb0 == opcode | 8'h90 == opcode | 8'h30 == opcode | 8'h10
     == opcode | 8'h50 == opcode | 8'h70 == opcode ? regs_sp : _GEN_1168; // @[CPU6502Core.scala 146:16 89:20]
  wire [15:0] _GEN_1188 = 8'hf0 == opcode | 8'hd0 == opcode | 8'hb0 == opcode | 8'h90 == opcode | 8'h30 == opcode | 8'h10
     == opcode | 8'h50 == opcode | 8'h70 == opcode ? execResult_result_newRegs_12_pc : _GEN_1169; // @[CPU6502Core.scala 146:16 89:20]
  wire  _GEN_1189 = 8'hf0 == opcode | 8'hd0 == opcode | 8'hb0 == opcode | 8'h90 == opcode | 8'h30 == opcode | 8'h10 ==
    opcode | 8'h50 == opcode | 8'h70 == opcode ? regs_flagC : _GEN_1170; // @[CPU6502Core.scala 146:16 89:20]
  wire  _GEN_1190 = 8'hf0 == opcode | 8'hd0 == opcode | 8'hb0 == opcode | 8'h90 == opcode | 8'h30 == opcode | 8'h10 ==
    opcode | 8'h50 == opcode | 8'h70 == opcode ? regs_flagZ : _GEN_1171; // @[CPU6502Core.scala 146:16 89:20]
  wire  _GEN_1191 = 8'hf0 == opcode | 8'hd0 == opcode | 8'hb0 == opcode | 8'h90 == opcode | 8'h30 == opcode | 8'h10 ==
    opcode | 8'h50 == opcode | 8'h70 == opcode ? regs_flagI : _GEN_1172; // @[CPU6502Core.scala 146:16 89:20]
  wire  _GEN_1192 = 8'hf0 == opcode | 8'hd0 == opcode | 8'hb0 == opcode | 8'h90 == opcode | 8'h30 == opcode | 8'h10 ==
    opcode | 8'h50 == opcode | 8'h70 == opcode ? regs_flagD : _GEN_1173; // @[CPU6502Core.scala 146:16 89:20]
  wire  _GEN_1194 = 8'hf0 == opcode | 8'hd0 == opcode | 8'hb0 == opcode | 8'h90 == opcode | 8'h30 == opcode | 8'h10 ==
    opcode | 8'h50 == opcode | 8'h70 == opcode ? regs_flagV : _GEN_1175; // @[CPU6502Core.scala 146:16 89:20]
  wire  _GEN_1195 = 8'hf0 == opcode | 8'hd0 == opcode | 8'hb0 == opcode | 8'h90 == opcode | 8'h30 == opcode | 8'h10 ==
    opcode | 8'h50 == opcode | 8'h70 == opcode ? regs_flagN : _GEN_1176; // @[CPU6502Core.scala 146:16 89:20]
  wire [15:0] _GEN_1196 = 8'hf0 == opcode | 8'hd0 == opcode | 8'hb0 == opcode | 8'h90 == opcode | 8'h30 == opcode | 8'h10
     == opcode | 8'h50 == opcode | 8'h70 == opcode ? regs_pc : _GEN_1177; // @[CPU6502Core.scala 146:16 89:20]
  wire [7:0] _GEN_1197 = 8'hf0 == opcode | 8'hd0 == opcode | 8'hb0 == opcode | 8'h90 == opcode | 8'h30 == opcode | 8'h10
     == opcode | 8'h50 == opcode | 8'h70 == opcode ? 8'h0 : _GEN_1178; // @[CPU6502Core.scala 146:16 89:20]
  wire  _GEN_1198 = 8'hf0 == opcode | 8'hd0 == opcode | 8'hb0 == opcode | 8'h90 == opcode | 8'h30 == opcode | 8'h10 ==
    opcode | 8'h50 == opcode | 8'h70 == opcode ? 1'h0 : _GEN_1179; // @[CPU6502Core.scala 146:16 89:20]
  wire  _GEN_1199 = 8'hf0 == opcode | 8'hd0 == opcode | 8'hb0 == opcode | 8'h90 == opcode | 8'h30 == opcode | 8'h10 ==
    opcode | 8'h50 == opcode | 8'h70 == opcode | _GEN_1180; // @[CPU6502Core.scala 146:16 89:20]
  wire [15:0] _GEN_1200 = 8'hf0 == opcode | 8'hd0 == opcode | 8'hb0 == opcode | 8'h90 == opcode | 8'h30 == opcode | 8'h10
     == opcode | 8'h50 == opcode | 8'h70 == opcode ? 16'h0 : _GEN_1181; // @[CPU6502Core.scala 146:16 89:20]
  wire  _GEN_1201 = 8'hc5 == opcode ? execResult_result_result_8_done : _GEN_1182; // @[CPU6502Core.scala 141:16 89:20]
  wire [2:0] _GEN_1202 = 8'hc5 == opcode ? execResult_result_result_8_nextCycle : _GEN_1183; // @[CPU6502Core.scala 141:16 89:20]
  wire [7:0] _GEN_1203 = 8'hc5 == opcode ? regs_a : _GEN_1184; // @[CPU6502Core.scala 141:16 89:20]
  wire [7:0] _GEN_1204 = 8'hc5 == opcode ? regs_x : _GEN_1185; // @[CPU6502Core.scala 141:16 89:20]
  wire [7:0] _GEN_1205 = 8'hc5 == opcode ? regs_y : _GEN_1186; // @[CPU6502Core.scala 141:16 89:20]
  wire [7:0] _GEN_1206 = 8'hc5 == opcode ? regs_sp : _GEN_1187; // @[CPU6502Core.scala 141:16 89:20]
  wire [15:0] _GEN_1207 = 8'hc5 == opcode ? execResult_result_newRegs_5_pc : _GEN_1188; // @[CPU6502Core.scala 141:16 89:20]
  wire  _GEN_1208 = 8'hc5 == opcode ? execResult_result_newRegs_11_flagC : _GEN_1189; // @[CPU6502Core.scala 141:16 89:20]
  wire  _GEN_1209 = 8'hc5 == opcode ? execResult_result_newRegs_11_flagZ : _GEN_1190; // @[CPU6502Core.scala 141:16 89:20]
  wire  _GEN_1210 = 8'hc5 == opcode ? regs_flagI : _GEN_1191; // @[CPU6502Core.scala 141:16 89:20]
  wire  _GEN_1211 = 8'hc5 == opcode ? regs_flagD : _GEN_1192; // @[CPU6502Core.scala 141:16 89:20]
  wire  _GEN_1213 = 8'hc5 == opcode ? regs_flagV : _GEN_1194; // @[CPU6502Core.scala 141:16 89:20]
  wire  _GEN_1214 = 8'hc5 == opcode ? execResult_result_newRegs_11_flagN : _GEN_1195; // @[CPU6502Core.scala 141:16 89:20]
  wire [15:0] _GEN_1215 = 8'hc5 == opcode ? execResult_result_result_8_memAddr : _GEN_1196; // @[CPU6502Core.scala 141:16 89:20]
  wire [7:0] _GEN_1216 = 8'hc5 == opcode ? 8'h0 : _GEN_1197; // @[CPU6502Core.scala 141:16 89:20]
  wire  _GEN_1217 = 8'hc5 == opcode ? 1'h0 : _GEN_1198; // @[CPU6502Core.scala 141:16 89:20]
  wire  _GEN_1218 = 8'hc5 == opcode ? execResult_result_result_6_memRead : _GEN_1199; // @[CPU6502Core.scala 141:16 89:20]
  wire [15:0] _GEN_1219 = 8'hc5 == opcode ? execResult_result_result_6_operand : _GEN_1200; // @[CPU6502Core.scala 141:16 89:20]
  wire  _GEN_1220 = 8'hc9 == opcode | 8'he0 == opcode | 8'hc0 == opcode | _GEN_1201; // @[CPU6502Core.scala 136:16 89:20]
  wire [2:0] _GEN_1221 = 8'hc9 == opcode | 8'he0 == opcode | 8'hc0 == opcode ? 3'h0 : _GEN_1202; // @[CPU6502Core.scala 136:16 89:20]
  wire [7:0] _GEN_1222 = 8'hc9 == opcode | 8'he0 == opcode | 8'hc0 == opcode ? regs_a : _GEN_1203; // @[CPU6502Core.scala 136:16 89:20]
  wire [7:0] _GEN_1223 = 8'hc9 == opcode | 8'he0 == opcode | 8'hc0 == opcode ? regs_x : _GEN_1204; // @[CPU6502Core.scala 136:16 89:20]
  wire [7:0] _GEN_1224 = 8'hc9 == opcode | 8'he0 == opcode | 8'hc0 == opcode ? regs_y : _GEN_1205; // @[CPU6502Core.scala 136:16 89:20]
  wire [7:0] _GEN_1225 = 8'hc9 == opcode | 8'he0 == opcode | 8'hc0 == opcode ? regs_sp : _GEN_1206; // @[CPU6502Core.scala 136:16 89:20]
  wire [15:0] _GEN_1226 = 8'hc9 == opcode | 8'he0 == opcode | 8'hc0 == opcode ? _regs_pc_T_1 : _GEN_1207; // @[CPU6502Core.scala 136:16 89:20]
  wire  _GEN_1227 = 8'hc9 == opcode | 8'he0 == opcode | 8'hc0 == opcode ? execResult_result_newRegs_10_flagC : _GEN_1208
    ; // @[CPU6502Core.scala 136:16 89:20]
  wire  _GEN_1228 = 8'hc9 == opcode | 8'he0 == opcode | 8'hc0 == opcode ? execResult_result_newRegs_10_flagZ : _GEN_1209
    ; // @[CPU6502Core.scala 136:16 89:20]
  wire  _GEN_1229 = 8'hc9 == opcode | 8'he0 == opcode | 8'hc0 == opcode ? regs_flagI : _GEN_1210; // @[CPU6502Core.scala 136:16 89:20]
  wire  _GEN_1230 = 8'hc9 == opcode | 8'he0 == opcode | 8'hc0 == opcode ? regs_flagD : _GEN_1211; // @[CPU6502Core.scala 136:16 89:20]
  wire  _GEN_1232 = 8'hc9 == opcode | 8'he0 == opcode | 8'hc0 == opcode ? regs_flagV : _GEN_1213; // @[CPU6502Core.scala 136:16 89:20]
  wire  _GEN_1233 = 8'hc9 == opcode | 8'he0 == opcode | 8'hc0 == opcode ? execResult_result_newRegs_10_flagN : _GEN_1214
    ; // @[CPU6502Core.scala 136:16 89:20]
  wire [15:0] _GEN_1234 = 8'hc9 == opcode | 8'he0 == opcode | 8'hc0 == opcode ? regs_pc : _GEN_1215; // @[CPU6502Core.scala 136:16 89:20]
  wire [7:0] _GEN_1235 = 8'hc9 == opcode | 8'he0 == opcode | 8'hc0 == opcode ? 8'h0 : _GEN_1216; // @[CPU6502Core.scala 136:16 89:20]
  wire  _GEN_1236 = 8'hc9 == opcode | 8'he0 == opcode | 8'hc0 == opcode ? 1'h0 : _GEN_1217; // @[CPU6502Core.scala 136:16 89:20]
  wire  _GEN_1237 = 8'hc9 == opcode | 8'he0 == opcode | 8'hc0 == opcode | _GEN_1218; // @[CPU6502Core.scala 136:16 89:20]
  wire [15:0] _GEN_1238 = 8'hc9 == opcode | 8'he0 == opcode | 8'hc0 == opcode ? 16'h0 : _GEN_1219; // @[CPU6502Core.scala 136:16 89:20]
  wire  _GEN_1239 = 8'h6 == opcode | 8'h46 == opcode | 8'h26 == opcode | 8'h66 == opcode ?
    execResult_result_result_6_done : _GEN_1220; // @[CPU6502Core.scala 131:16 89:20]
  wire [2:0] _GEN_1240 = 8'h6 == opcode | 8'h46 == opcode | 8'h26 == opcode | 8'h66 == opcode ?
    execResult_result_result_6_nextCycle : _GEN_1221; // @[CPU6502Core.scala 131:16 89:20]
  wire [7:0] _GEN_1241 = 8'h6 == opcode | 8'h46 == opcode | 8'h26 == opcode | 8'h66 == opcode ? regs_a : _GEN_1222; // @[CPU6502Core.scala 131:16 89:20]
  wire [7:0] _GEN_1242 = 8'h6 == opcode | 8'h46 == opcode | 8'h26 == opcode | 8'h66 == opcode ? regs_x : _GEN_1223; // @[CPU6502Core.scala 131:16 89:20]
  wire [7:0] _GEN_1243 = 8'h6 == opcode | 8'h46 == opcode | 8'h26 == opcode | 8'h66 == opcode ? regs_y : _GEN_1224; // @[CPU6502Core.scala 131:16 89:20]
  wire [7:0] _GEN_1244 = 8'h6 == opcode | 8'h46 == opcode | 8'h26 == opcode | 8'h66 == opcode ? regs_sp : _GEN_1225; // @[CPU6502Core.scala 131:16 89:20]
  wire [15:0] _GEN_1245 = 8'h6 == opcode | 8'h46 == opcode | 8'h26 == opcode | 8'h66 == opcode ?
    execResult_result_newRegs_5_pc : _GEN_1226; // @[CPU6502Core.scala 131:16 89:20]
  wire  _GEN_1246 = 8'h6 == opcode | 8'h46 == opcode | 8'h26 == opcode | 8'h66 == opcode ?
    execResult_result_newRegs_9_flagC : _GEN_1227; // @[CPU6502Core.scala 131:16 89:20]
  wire  _GEN_1247 = 8'h6 == opcode | 8'h46 == opcode | 8'h26 == opcode | 8'h66 == opcode ?
    execResult_result_newRegs_9_flagZ : _GEN_1228; // @[CPU6502Core.scala 131:16 89:20]
  wire  _GEN_1248 = 8'h6 == opcode | 8'h46 == opcode | 8'h26 == opcode | 8'h66 == opcode ? regs_flagI : _GEN_1229; // @[CPU6502Core.scala 131:16 89:20]
  wire  _GEN_1249 = 8'h6 == opcode | 8'h46 == opcode | 8'h26 == opcode | 8'h66 == opcode ? regs_flagD : _GEN_1230; // @[CPU6502Core.scala 131:16 89:20]
  wire  _GEN_1251 = 8'h6 == opcode | 8'h46 == opcode | 8'h26 == opcode | 8'h66 == opcode ? regs_flagV : _GEN_1232; // @[CPU6502Core.scala 131:16 89:20]
  wire  _GEN_1252 = 8'h6 == opcode | 8'h46 == opcode | 8'h26 == opcode | 8'h66 == opcode ?
    execResult_result_newRegs_9_flagN : _GEN_1233; // @[CPU6502Core.scala 131:16 89:20]
  wire [15:0] _GEN_1253 = 8'h6 == opcode | 8'h46 == opcode | 8'h26 == opcode | 8'h66 == opcode ?
    execResult_result_result_6_memAddr : _GEN_1234; // @[CPU6502Core.scala 131:16 89:20]
  wire [7:0] _GEN_1254 = 8'h6 == opcode | 8'h46 == opcode | 8'h26 == opcode | 8'h66 == opcode ?
    execResult_result_result_10_memData : _GEN_1235; // @[CPU6502Core.scala 131:16 89:20]
  wire  _GEN_1255 = 8'h6 == opcode | 8'h46 == opcode | 8'h26 == opcode | 8'h66 == opcode ?
    execResult_result_result_6_done : _GEN_1236; // @[CPU6502Core.scala 131:16 89:20]
  wire  _GEN_1256 = 8'h6 == opcode | 8'h46 == opcode | 8'h26 == opcode | 8'h66 == opcode ?
    execResult_result_result_6_memRead : _GEN_1237; // @[CPU6502Core.scala 131:16 89:20]
  wire [15:0] _GEN_1257 = 8'h6 == opcode | 8'h46 == opcode | 8'h26 == opcode | 8'h66 == opcode ?
    execResult_result_result_6_operand : _GEN_1238; // @[CPU6502Core.scala 131:16 89:20]
  wire  _GEN_1258 = 8'ha == opcode | 8'h4a == opcode | 8'h2a == opcode | 8'h6a == opcode | _GEN_1239; // @[CPU6502Core.scala 126:16 89:20]
  wire [2:0] _GEN_1259 = 8'ha == opcode | 8'h4a == opcode | 8'h2a == opcode | 8'h6a == opcode ? 3'h0 : _GEN_1240; // @[CPU6502Core.scala 126:16 89:20]
  wire [7:0] _GEN_1260 = 8'ha == opcode | 8'h4a == opcode | 8'h2a == opcode | 8'h6a == opcode ? execResult_result_res_8
     : _GEN_1241; // @[CPU6502Core.scala 126:16 89:20]
  wire [7:0] _GEN_1261 = 8'ha == opcode | 8'h4a == opcode | 8'h2a == opcode | 8'h6a == opcode ? regs_x : _GEN_1242; // @[CPU6502Core.scala 126:16 89:20]
  wire [7:0] _GEN_1262 = 8'ha == opcode | 8'h4a == opcode | 8'h2a == opcode | 8'h6a == opcode ? regs_y : _GEN_1243; // @[CPU6502Core.scala 126:16 89:20]
  wire [7:0] _GEN_1263 = 8'ha == opcode | 8'h4a == opcode | 8'h2a == opcode | 8'h6a == opcode ? regs_sp : _GEN_1244; // @[CPU6502Core.scala 126:16 89:20]
  wire [15:0] _GEN_1264 = 8'ha == opcode | 8'h4a == opcode | 8'h2a == opcode | 8'h6a == opcode ? regs_pc : _GEN_1245; // @[CPU6502Core.scala 126:16 89:20]
  wire  _GEN_1265 = 8'ha == opcode | 8'h4a == opcode | 8'h2a == opcode | 8'h6a == opcode ?
    execResult_result_newRegs_8_flagC : _GEN_1246; // @[CPU6502Core.scala 126:16 89:20]
  wire  _GEN_1266 = 8'ha == opcode | 8'h4a == opcode | 8'h2a == opcode | 8'h6a == opcode ?
    execResult_result_newRegs_8_flagZ : _GEN_1247; // @[CPU6502Core.scala 126:16 89:20]
  wire  _GEN_1267 = 8'ha == opcode | 8'h4a == opcode | 8'h2a == opcode | 8'h6a == opcode ? regs_flagI : _GEN_1248; // @[CPU6502Core.scala 126:16 89:20]
  wire  _GEN_1268 = 8'ha == opcode | 8'h4a == opcode | 8'h2a == opcode | 8'h6a == opcode ? regs_flagD : _GEN_1249; // @[CPU6502Core.scala 126:16 89:20]
  wire  _GEN_1270 = 8'ha == opcode | 8'h4a == opcode | 8'h2a == opcode | 8'h6a == opcode ? regs_flagV : _GEN_1251; // @[CPU6502Core.scala 126:16 89:20]
  wire  _GEN_1271 = 8'ha == opcode | 8'h4a == opcode | 8'h2a == opcode | 8'h6a == opcode ?
    execResult_result_newRegs_8_flagN : _GEN_1252; // @[CPU6502Core.scala 126:16 89:20]
  wire [15:0] _GEN_1272 = 8'ha == opcode | 8'h4a == opcode | 8'h2a == opcode | 8'h6a == opcode ? 16'h0 : _GEN_1253; // @[CPU6502Core.scala 126:16 89:20]
  wire [7:0] _GEN_1273 = 8'ha == opcode | 8'h4a == opcode | 8'h2a == opcode | 8'h6a == opcode ? 8'h0 : _GEN_1254; // @[CPU6502Core.scala 126:16 89:20]
  wire  _GEN_1274 = 8'ha == opcode | 8'h4a == opcode | 8'h2a == opcode | 8'h6a == opcode ? 1'h0 : _GEN_1255; // @[CPU6502Core.scala 126:16 89:20]
  wire  _GEN_1275 = 8'ha == opcode | 8'h4a == opcode | 8'h2a == opcode | 8'h6a == opcode ? 1'h0 : _GEN_1256; // @[CPU6502Core.scala 126:16 89:20]
  wire [15:0] _GEN_1276 = 8'ha == opcode | 8'h4a == opcode | 8'h2a == opcode | 8'h6a == opcode ? 16'h0 : _GEN_1257; // @[CPU6502Core.scala 126:16 89:20]
  wire  _GEN_1277 = 8'h24 == opcode ? execResult_result_result_8_done : _GEN_1258; // @[CPU6502Core.scala 121:16 89:20]
  wire [2:0] _GEN_1278 = 8'h24 == opcode ? execResult_result_result_8_nextCycle : _GEN_1259; // @[CPU6502Core.scala 121:16 89:20]
  wire [7:0] _GEN_1279 = 8'h24 == opcode ? regs_a : _GEN_1260; // @[CPU6502Core.scala 121:16 89:20]
  wire [7:0] _GEN_1280 = 8'h24 == opcode ? regs_x : _GEN_1261; // @[CPU6502Core.scala 121:16 89:20]
  wire [7:0] _GEN_1281 = 8'h24 == opcode ? regs_y : _GEN_1262; // @[CPU6502Core.scala 121:16 89:20]
  wire [7:0] _GEN_1282 = 8'h24 == opcode ? regs_sp : _GEN_1263; // @[CPU6502Core.scala 121:16 89:20]
  wire [15:0] _GEN_1283 = 8'h24 == opcode ? execResult_result_newRegs_5_pc : _GEN_1264; // @[CPU6502Core.scala 121:16 89:20]
  wire  _GEN_1284 = 8'h24 == opcode ? regs_flagC : _GEN_1265; // @[CPU6502Core.scala 121:16 89:20]
  wire  _GEN_1285 = 8'h24 == opcode ? execResult_result_newRegs_7_flagZ : _GEN_1266; // @[CPU6502Core.scala 121:16 89:20]
  wire  _GEN_1286 = 8'h24 == opcode ? regs_flagI : _GEN_1267; // @[CPU6502Core.scala 121:16 89:20]
  wire  _GEN_1287 = 8'h24 == opcode ? regs_flagD : _GEN_1268; // @[CPU6502Core.scala 121:16 89:20]
  wire  _GEN_1289 = 8'h24 == opcode ? execResult_result_newRegs_7_flagV : _GEN_1270; // @[CPU6502Core.scala 121:16 89:20]
  wire  _GEN_1290 = 8'h24 == opcode ? execResult_result_newRegs_7_flagN : _GEN_1271; // @[CPU6502Core.scala 121:16 89:20]
  wire [15:0] _GEN_1291 = 8'h24 == opcode ? execResult_result_result_8_memAddr : _GEN_1272; // @[CPU6502Core.scala 121:16 89:20]
  wire [7:0] _GEN_1292 = 8'h24 == opcode ? 8'h0 : _GEN_1273; // @[CPU6502Core.scala 121:16 89:20]
  wire  _GEN_1293 = 8'h24 == opcode ? 1'h0 : _GEN_1274; // @[CPU6502Core.scala 121:16 89:20]
  wire  _GEN_1294 = 8'h24 == opcode ? execResult_result_result_6_memRead : _GEN_1275; // @[CPU6502Core.scala 121:16 89:20]
  wire [15:0] _GEN_1295 = 8'h24 == opcode ? execResult_result_result_6_operand : _GEN_1276; // @[CPU6502Core.scala 121:16 89:20]
  wire  _GEN_1296 = 8'h29 == opcode | 8'h9 == opcode | 8'h49 == opcode | _GEN_1277; // @[CPU6502Core.scala 116:16 89:20]
  wire [2:0] _GEN_1297 = 8'h29 == opcode | 8'h9 == opcode | 8'h49 == opcode ? 3'h0 : _GEN_1278; // @[CPU6502Core.scala 116:16 89:20]
  wire [7:0] _GEN_1298 = 8'h29 == opcode | 8'h9 == opcode | 8'h49 == opcode ? execResult_result_res_7 : _GEN_1279; // @[CPU6502Core.scala 116:16 89:20]
  wire [7:0] _GEN_1299 = 8'h29 == opcode | 8'h9 == opcode | 8'h49 == opcode ? regs_x : _GEN_1280; // @[CPU6502Core.scala 116:16 89:20]
  wire [7:0] _GEN_1300 = 8'h29 == opcode | 8'h9 == opcode | 8'h49 == opcode ? regs_y : _GEN_1281; // @[CPU6502Core.scala 116:16 89:20]
  wire [7:0] _GEN_1301 = 8'h29 == opcode | 8'h9 == opcode | 8'h49 == opcode ? regs_sp : _GEN_1282; // @[CPU6502Core.scala 116:16 89:20]
  wire [15:0] _GEN_1302 = 8'h29 == opcode | 8'h9 == opcode | 8'h49 == opcode ? _regs_pc_T_1 : _GEN_1283; // @[CPU6502Core.scala 116:16 89:20]
  wire  _GEN_1303 = 8'h29 == opcode | 8'h9 == opcode | 8'h49 == opcode ? regs_flagC : _GEN_1284; // @[CPU6502Core.scala 116:16 89:20]
  wire  _GEN_1304 = 8'h29 == opcode | 8'h9 == opcode | 8'h49 == opcode ? execResult_result_newRegs_6_flagZ : _GEN_1285; // @[CPU6502Core.scala 116:16 89:20]
  wire  _GEN_1305 = 8'h29 == opcode | 8'h9 == opcode | 8'h49 == opcode ? regs_flagI : _GEN_1286; // @[CPU6502Core.scala 116:16 89:20]
  wire  _GEN_1306 = 8'h29 == opcode | 8'h9 == opcode | 8'h49 == opcode ? regs_flagD : _GEN_1287; // @[CPU6502Core.scala 116:16 89:20]
  wire  _GEN_1308 = 8'h29 == opcode | 8'h9 == opcode | 8'h49 == opcode ? regs_flagV : _GEN_1289; // @[CPU6502Core.scala 116:16 89:20]
  wire  _GEN_1309 = 8'h29 == opcode | 8'h9 == opcode | 8'h49 == opcode ? execResult_result_newRegs_6_flagN : _GEN_1290; // @[CPU6502Core.scala 116:16 89:20]
  wire [15:0] _GEN_1310 = 8'h29 == opcode | 8'h9 == opcode | 8'h49 == opcode ? regs_pc : _GEN_1291; // @[CPU6502Core.scala 116:16 89:20]
  wire [7:0] _GEN_1311 = 8'h29 == opcode | 8'h9 == opcode | 8'h49 == opcode ? 8'h0 : _GEN_1292; // @[CPU6502Core.scala 116:16 89:20]
  wire  _GEN_1312 = 8'h29 == opcode | 8'h9 == opcode | 8'h49 == opcode ? 1'h0 : _GEN_1293; // @[CPU6502Core.scala 116:16 89:20]
  wire  _GEN_1313 = 8'h29 == opcode | 8'h9 == opcode | 8'h49 == opcode | _GEN_1294; // @[CPU6502Core.scala 116:16 89:20]
  wire [15:0] _GEN_1314 = 8'h29 == opcode | 8'h9 == opcode | 8'h49 == opcode ? 16'h0 : _GEN_1295; // @[CPU6502Core.scala 116:16 89:20]
  wire  _GEN_1315 = 8'he6 == opcode | 8'hc6 == opcode ? execResult_result_result_6_done : _GEN_1296; // @[CPU6502Core.scala 111:16 89:20]
  wire [2:0] _GEN_1316 = 8'he6 == opcode | 8'hc6 == opcode ? execResult_result_result_6_nextCycle : _GEN_1297; // @[CPU6502Core.scala 111:16 89:20]
  wire [7:0] _GEN_1317 = 8'he6 == opcode | 8'hc6 == opcode ? regs_a : _GEN_1298; // @[CPU6502Core.scala 111:16 89:20]
  wire [7:0] _GEN_1318 = 8'he6 == opcode | 8'hc6 == opcode ? regs_x : _GEN_1299; // @[CPU6502Core.scala 111:16 89:20]
  wire [7:0] _GEN_1319 = 8'he6 == opcode | 8'hc6 == opcode ? regs_y : _GEN_1300; // @[CPU6502Core.scala 111:16 89:20]
  wire [7:0] _GEN_1320 = 8'he6 == opcode | 8'hc6 == opcode ? regs_sp : _GEN_1301; // @[CPU6502Core.scala 111:16 89:20]
  wire [15:0] _GEN_1321 = 8'he6 == opcode | 8'hc6 == opcode ? execResult_result_newRegs_5_pc : _GEN_1302; // @[CPU6502Core.scala 111:16 89:20]
  wire  _GEN_1322 = 8'he6 == opcode | 8'hc6 == opcode ? regs_flagC : _GEN_1303; // @[CPU6502Core.scala 111:16 89:20]
  wire  _GEN_1323 = 8'he6 == opcode | 8'hc6 == opcode ? execResult_result_newRegs_5_flagZ : _GEN_1304; // @[CPU6502Core.scala 111:16 89:20]
  wire  _GEN_1324 = 8'he6 == opcode | 8'hc6 == opcode ? regs_flagI : _GEN_1305; // @[CPU6502Core.scala 111:16 89:20]
  wire  _GEN_1325 = 8'he6 == opcode | 8'hc6 == opcode ? regs_flagD : _GEN_1306; // @[CPU6502Core.scala 111:16 89:20]
  wire  _GEN_1327 = 8'he6 == opcode | 8'hc6 == opcode ? regs_flagV : _GEN_1308; // @[CPU6502Core.scala 111:16 89:20]
  wire  _GEN_1328 = 8'he6 == opcode | 8'hc6 == opcode ? execResult_result_newRegs_5_flagN : _GEN_1309; // @[CPU6502Core.scala 111:16 89:20]
  wire [15:0] _GEN_1329 = 8'he6 == opcode | 8'hc6 == opcode ? execResult_result_result_6_memAddr : _GEN_1310; // @[CPU6502Core.scala 111:16 89:20]
  wire [7:0] _GEN_1330 = 8'he6 == opcode | 8'hc6 == opcode ? execResult_result_result_6_memData : _GEN_1311; // @[CPU6502Core.scala 111:16 89:20]
  wire  _GEN_1331 = 8'he6 == opcode | 8'hc6 == opcode ? execResult_result_result_6_done : _GEN_1312; // @[CPU6502Core.scala 111:16 89:20]
  wire  _GEN_1332 = 8'he6 == opcode | 8'hc6 == opcode ? execResult_result_result_6_memRead : _GEN_1313; // @[CPU6502Core.scala 111:16 89:20]
  wire [15:0] _GEN_1333 = 8'he6 == opcode | 8'hc6 == opcode ? execResult_result_result_6_operand : _GEN_1314; // @[CPU6502Core.scala 111:16 89:20]
  wire  _GEN_1334 = 8'he9 == opcode | _GEN_1315; // @[CPU6502Core.scala 89:20 107:27]
  wire [2:0] _GEN_1335 = 8'he9 == opcode ? 3'h0 : _GEN_1316; // @[CPU6502Core.scala 89:20 107:27]
  wire [7:0] _GEN_1336 = 8'he9 == opcode ? execResult_result_newRegs_4_a : _GEN_1317; // @[CPU6502Core.scala 89:20 107:27]
  wire [7:0] _GEN_1337 = 8'he9 == opcode ? regs_x : _GEN_1318; // @[CPU6502Core.scala 89:20 107:27]
  wire [7:0] _GEN_1338 = 8'he9 == opcode ? regs_y : _GEN_1319; // @[CPU6502Core.scala 89:20 107:27]
  wire [7:0] _GEN_1339 = 8'he9 == opcode ? regs_sp : _GEN_1320; // @[CPU6502Core.scala 89:20 107:27]
  wire [15:0] _GEN_1340 = 8'he9 == opcode ? _regs_pc_T_1 : _GEN_1321; // @[CPU6502Core.scala 89:20 107:27]
  wire  _GEN_1341 = 8'he9 == opcode ? execResult_result_newRegs_4_flagC : _GEN_1322; // @[CPU6502Core.scala 89:20 107:27]
  wire  _GEN_1342 = 8'he9 == opcode ? execResult_result_newRegs_4_flagZ : _GEN_1323; // @[CPU6502Core.scala 89:20 107:27]
  wire  _GEN_1343 = 8'he9 == opcode ? regs_flagI : _GEN_1324; // @[CPU6502Core.scala 89:20 107:27]
  wire  _GEN_1344 = 8'he9 == opcode ? regs_flagD : _GEN_1325; // @[CPU6502Core.scala 89:20 107:27]
  wire  _GEN_1346 = 8'he9 == opcode ? execResult_result_newRegs_4_flagV : _GEN_1327; // @[CPU6502Core.scala 89:20 107:27]
  wire  _GEN_1347 = 8'he9 == opcode ? execResult_result_newRegs_4_flagN : _GEN_1328; // @[CPU6502Core.scala 89:20 107:27]
  wire [15:0] _GEN_1348 = 8'he9 == opcode ? regs_pc : _GEN_1329; // @[CPU6502Core.scala 89:20 107:27]
  wire [7:0] _GEN_1349 = 8'he9 == opcode ? 8'h0 : _GEN_1330; // @[CPU6502Core.scala 89:20 107:27]
  wire  _GEN_1350 = 8'he9 == opcode ? 1'h0 : _GEN_1331; // @[CPU6502Core.scala 89:20 107:27]
  wire  _GEN_1351 = 8'he9 == opcode | _GEN_1332; // @[CPU6502Core.scala 89:20 107:27]
  wire [15:0] _GEN_1352 = 8'he9 == opcode ? 16'h0 : _GEN_1333; // @[CPU6502Core.scala 89:20 107:27]
  wire  _GEN_1353 = 8'h69 == opcode | _GEN_1334; // @[CPU6502Core.scala 89:20 106:27]
  wire [2:0] _GEN_1354 = 8'h69 == opcode ? 3'h0 : _GEN_1335; // @[CPU6502Core.scala 89:20 106:27]
  wire [7:0] _GEN_1355 = 8'h69 == opcode ? execResult_result_newRegs_3_a : _GEN_1336; // @[CPU6502Core.scala 89:20 106:27]
  wire [7:0] _GEN_1356 = 8'h69 == opcode ? regs_x : _GEN_1337; // @[CPU6502Core.scala 89:20 106:27]
  wire [7:0] _GEN_1357 = 8'h69 == opcode ? regs_y : _GEN_1338; // @[CPU6502Core.scala 89:20 106:27]
  wire [7:0] _GEN_1358 = 8'h69 == opcode ? regs_sp : _GEN_1339; // @[CPU6502Core.scala 89:20 106:27]
  wire [15:0] _GEN_1359 = 8'h69 == opcode ? _regs_pc_T_1 : _GEN_1340; // @[CPU6502Core.scala 89:20 106:27]
  wire  _GEN_1360 = 8'h69 == opcode ? execResult_result_newRegs_3_flagC : _GEN_1341; // @[CPU6502Core.scala 89:20 106:27]
  wire  _GEN_1361 = 8'h69 == opcode ? execResult_result_newRegs_3_flagZ : _GEN_1342; // @[CPU6502Core.scala 89:20 106:27]
  wire  _GEN_1362 = 8'h69 == opcode ? regs_flagI : _GEN_1343; // @[CPU6502Core.scala 89:20 106:27]
  wire  _GEN_1363 = 8'h69 == opcode ? regs_flagD : _GEN_1344; // @[CPU6502Core.scala 89:20 106:27]
  wire  _GEN_1365 = 8'h69 == opcode ? execResult_result_newRegs_3_flagV : _GEN_1346; // @[CPU6502Core.scala 89:20 106:27]
  wire  _GEN_1366 = 8'h69 == opcode ? execResult_result_newRegs_3_flagN : _GEN_1347; // @[CPU6502Core.scala 89:20 106:27]
  wire [15:0] _GEN_1367 = 8'h69 == opcode ? regs_pc : _GEN_1348; // @[CPU6502Core.scala 89:20 106:27]
  wire [7:0] _GEN_1368 = 8'h69 == opcode ? 8'h0 : _GEN_1349; // @[CPU6502Core.scala 89:20 106:27]
  wire  _GEN_1369 = 8'h69 == opcode ? 1'h0 : _GEN_1350; // @[CPU6502Core.scala 89:20 106:27]
  wire  _GEN_1370 = 8'h69 == opcode | _GEN_1351; // @[CPU6502Core.scala 89:20 106:27]
  wire [15:0] _GEN_1371 = 8'h69 == opcode ? 16'h0 : _GEN_1352; // @[CPU6502Core.scala 89:20 106:27]
  wire  _GEN_1372 = 8'he8 == opcode | 8'hc8 == opcode | 8'hca == opcode | 8'h88 == opcode | 8'h1a == opcode | 8'h3a ==
    opcode | _GEN_1353; // @[CPU6502Core.scala 102:16 89:20]
  wire [2:0] _GEN_1373 = 8'he8 == opcode | 8'hc8 == opcode | 8'hca == opcode | 8'h88 == opcode | 8'h1a == opcode | 8'h3a
     == opcode ? 3'h0 : _GEN_1354; // @[CPU6502Core.scala 102:16 89:20]
  wire [7:0] _GEN_1374 = 8'he8 == opcode | 8'hc8 == opcode | 8'hca == opcode | 8'h88 == opcode | 8'h1a == opcode | 8'h3a
     == opcode ? execResult_result_newRegs_2_a : _GEN_1355; // @[CPU6502Core.scala 102:16 89:20]
  wire [7:0] _GEN_1375 = 8'he8 == opcode | 8'hc8 == opcode | 8'hca == opcode | 8'h88 == opcode | 8'h1a == opcode | 8'h3a
     == opcode ? execResult_result_newRegs_2_x : _GEN_1356; // @[CPU6502Core.scala 102:16 89:20]
  wire [7:0] _GEN_1376 = 8'he8 == opcode | 8'hc8 == opcode | 8'hca == opcode | 8'h88 == opcode | 8'h1a == opcode | 8'h3a
     == opcode ? execResult_result_newRegs_2_y : _GEN_1357; // @[CPU6502Core.scala 102:16 89:20]
  wire [7:0] _GEN_1377 = 8'he8 == opcode | 8'hc8 == opcode | 8'hca == opcode | 8'h88 == opcode | 8'h1a == opcode | 8'h3a
     == opcode ? regs_sp : _GEN_1358; // @[CPU6502Core.scala 102:16 89:20]
  wire [15:0] _GEN_1378 = 8'he8 == opcode | 8'hc8 == opcode | 8'hca == opcode | 8'h88 == opcode | 8'h1a == opcode | 8'h3a
     == opcode ? regs_pc : _GEN_1359; // @[CPU6502Core.scala 102:16 89:20]
  wire  _GEN_1379 = 8'he8 == opcode | 8'hc8 == opcode | 8'hca == opcode | 8'h88 == opcode | 8'h1a == opcode | 8'h3a ==
    opcode ? regs_flagC : _GEN_1360; // @[CPU6502Core.scala 102:16 89:20]
  wire  _GEN_1380 = 8'he8 == opcode | 8'hc8 == opcode | 8'hca == opcode | 8'h88 == opcode | 8'h1a == opcode | 8'h3a ==
    opcode ? execResult_result_newRegs_2_flagZ : _GEN_1361; // @[CPU6502Core.scala 102:16 89:20]
  wire  _GEN_1381 = 8'he8 == opcode | 8'hc8 == opcode | 8'hca == opcode | 8'h88 == opcode | 8'h1a == opcode | 8'h3a ==
    opcode ? regs_flagI : _GEN_1362; // @[CPU6502Core.scala 102:16 89:20]
  wire  _GEN_1382 = 8'he8 == opcode | 8'hc8 == opcode | 8'hca == opcode | 8'h88 == opcode | 8'h1a == opcode | 8'h3a ==
    opcode ? regs_flagD : _GEN_1363; // @[CPU6502Core.scala 102:16 89:20]
  wire  _GEN_1384 = 8'he8 == opcode | 8'hc8 == opcode | 8'hca == opcode | 8'h88 == opcode | 8'h1a == opcode | 8'h3a ==
    opcode ? regs_flagV : _GEN_1365; // @[CPU6502Core.scala 102:16 89:20]
  wire  _GEN_1385 = 8'he8 == opcode | 8'hc8 == opcode | 8'hca == opcode | 8'h88 == opcode | 8'h1a == opcode | 8'h3a ==
    opcode ? execResult_result_newRegs_2_flagN : _GEN_1366; // @[CPU6502Core.scala 102:16 89:20]
  wire [15:0] _GEN_1386 = 8'he8 == opcode | 8'hc8 == opcode | 8'hca == opcode | 8'h88 == opcode | 8'h1a == opcode | 8'h3a
     == opcode ? 16'h0 : _GEN_1367; // @[CPU6502Core.scala 102:16 89:20]
  wire [7:0] _GEN_1387 = 8'he8 == opcode | 8'hc8 == opcode | 8'hca == opcode | 8'h88 == opcode | 8'h1a == opcode | 8'h3a
     == opcode ? 8'h0 : _GEN_1368; // @[CPU6502Core.scala 102:16 89:20]
  wire  _GEN_1388 = 8'he8 == opcode | 8'hc8 == opcode | 8'hca == opcode | 8'h88 == opcode | 8'h1a == opcode | 8'h3a ==
    opcode ? 1'h0 : _GEN_1369; // @[CPU6502Core.scala 102:16 89:20]
  wire  _GEN_1389 = 8'he8 == opcode | 8'hc8 == opcode | 8'hca == opcode | 8'h88 == opcode | 8'h1a == opcode | 8'h3a ==
    opcode ? 1'h0 : _GEN_1370; // @[CPU6502Core.scala 102:16 89:20]
  wire [15:0] _GEN_1390 = 8'he8 == opcode | 8'hc8 == opcode | 8'hca == opcode | 8'h88 == opcode | 8'h1a == opcode | 8'h3a
     == opcode ? 16'h0 : _GEN_1371; // @[CPU6502Core.scala 102:16 89:20]
  wire  _GEN_1391 = 8'haa == opcode | 8'ha8 == opcode | 8'h8a == opcode | 8'h98 == opcode | 8'hba == opcode | 8'h9a ==
    opcode | _GEN_1372; // @[CPU6502Core.scala 89:20 97:16]
  wire [2:0] _GEN_1392 = 8'haa == opcode | 8'ha8 == opcode | 8'h8a == opcode | 8'h98 == opcode | 8'hba == opcode | 8'h9a
     == opcode ? 3'h0 : _GEN_1373; // @[CPU6502Core.scala 89:20 97:16]
  wire [7:0] _GEN_1393 = 8'haa == opcode | 8'ha8 == opcode | 8'h8a == opcode | 8'h98 == opcode | 8'hba == opcode | 8'h9a
     == opcode ? execResult_result_newRegs_1_a : _GEN_1374; // @[CPU6502Core.scala 89:20 97:16]
  wire [7:0] _GEN_1394 = 8'haa == opcode | 8'ha8 == opcode | 8'h8a == opcode | 8'h98 == opcode | 8'hba == opcode | 8'h9a
     == opcode ? execResult_result_newRegs_1_x : _GEN_1375; // @[CPU6502Core.scala 89:20 97:16]
  wire [7:0] _GEN_1395 = 8'haa == opcode | 8'ha8 == opcode | 8'h8a == opcode | 8'h98 == opcode | 8'hba == opcode | 8'h9a
     == opcode ? execResult_result_newRegs_1_y : _GEN_1376; // @[CPU6502Core.scala 89:20 97:16]
  wire [7:0] _GEN_1396 = 8'haa == opcode | 8'ha8 == opcode | 8'h8a == opcode | 8'h98 == opcode | 8'hba == opcode | 8'h9a
     == opcode ? execResult_result_newRegs_1_sp : _GEN_1377; // @[CPU6502Core.scala 89:20 97:16]
  wire [15:0] _GEN_1397 = 8'haa == opcode | 8'ha8 == opcode | 8'h8a == opcode | 8'h98 == opcode | 8'hba == opcode | 8'h9a
     == opcode ? regs_pc : _GEN_1378; // @[CPU6502Core.scala 89:20 97:16]
  wire  _GEN_1398 = 8'haa == opcode | 8'ha8 == opcode | 8'h8a == opcode | 8'h98 == opcode | 8'hba == opcode | 8'h9a ==
    opcode ? regs_flagC : _GEN_1379; // @[CPU6502Core.scala 89:20 97:16]
  wire  _GEN_1399 = 8'haa == opcode | 8'ha8 == opcode | 8'h8a == opcode | 8'h98 == opcode | 8'hba == opcode | 8'h9a ==
    opcode ? execResult_result_newRegs_1_flagZ : _GEN_1380; // @[CPU6502Core.scala 89:20 97:16]
  wire  _GEN_1400 = 8'haa == opcode | 8'ha8 == opcode | 8'h8a == opcode | 8'h98 == opcode | 8'hba == opcode | 8'h9a ==
    opcode ? regs_flagI : _GEN_1381; // @[CPU6502Core.scala 89:20 97:16]
  wire  _GEN_1401 = 8'haa == opcode | 8'ha8 == opcode | 8'h8a == opcode | 8'h98 == opcode | 8'hba == opcode | 8'h9a ==
    opcode ? regs_flagD : _GEN_1382; // @[CPU6502Core.scala 89:20 97:16]
  wire  _GEN_1403 = 8'haa == opcode | 8'ha8 == opcode | 8'h8a == opcode | 8'h98 == opcode | 8'hba == opcode | 8'h9a ==
    opcode ? regs_flagV : _GEN_1384; // @[CPU6502Core.scala 89:20 97:16]
  wire  _GEN_1404 = 8'haa == opcode | 8'ha8 == opcode | 8'h8a == opcode | 8'h98 == opcode | 8'hba == opcode | 8'h9a ==
    opcode ? execResult_result_newRegs_1_flagN : _GEN_1385; // @[CPU6502Core.scala 89:20 97:16]
  wire [15:0] _GEN_1405 = 8'haa == opcode | 8'ha8 == opcode | 8'h8a == opcode | 8'h98 == opcode | 8'hba == opcode | 8'h9a
     == opcode ? 16'h0 : _GEN_1386; // @[CPU6502Core.scala 89:20 97:16]
  wire [7:0] _GEN_1406 = 8'haa == opcode | 8'ha8 == opcode | 8'h8a == opcode | 8'h98 == opcode | 8'hba == opcode | 8'h9a
     == opcode ? 8'h0 : _GEN_1387; // @[CPU6502Core.scala 89:20 97:16]
  wire  _GEN_1407 = 8'haa == opcode | 8'ha8 == opcode | 8'h8a == opcode | 8'h98 == opcode | 8'hba == opcode | 8'h9a ==
    opcode ? 1'h0 : _GEN_1388; // @[CPU6502Core.scala 89:20 97:16]
  wire  _GEN_1408 = 8'haa == opcode | 8'ha8 == opcode | 8'h8a == opcode | 8'h98 == opcode | 8'hba == opcode | 8'h9a ==
    opcode ? 1'h0 : _GEN_1389; // @[CPU6502Core.scala 89:20 97:16]
  wire [15:0] _GEN_1409 = 8'haa == opcode | 8'ha8 == opcode | 8'h8a == opcode | 8'h98 == opcode | 8'hba == opcode | 8'h9a
     == opcode ? 16'h0 : _GEN_1390; // @[CPU6502Core.scala 89:20 97:16]
  wire  execResult_result_1_done = 8'h18 == opcode | 8'h38 == opcode | 8'hd8 == opcode | 8'hf8 == opcode | 8'h58 ==
    opcode | 8'h78 == opcode | 8'hb8 == opcode | 8'hea == opcode | _GEN_1391; // @[CPU6502Core.scala 89:20 92:16]
  wire [2:0] execResult_result_1_nextCycle = 8'h18 == opcode | 8'h38 == opcode | 8'hd8 == opcode | 8'hf8 == opcode | 8'h58
     == opcode | 8'h78 == opcode | 8'hb8 == opcode | 8'hea == opcode ? 3'h0 : _GEN_1392; // @[CPU6502Core.scala 89:20 92:16]
  wire [7:0] execResult_result_1_regs_a = 8'h18 == opcode | 8'h38 == opcode | 8'hd8 == opcode | 8'hf8 == opcode | 8'h58
     == opcode | 8'h78 == opcode | 8'hb8 == opcode | 8'hea == opcode ? regs_a : _GEN_1393; // @[CPU6502Core.scala 89:20 92:16]
  wire [7:0] execResult_result_1_regs_x = 8'h18 == opcode | 8'h38 == opcode | 8'hd8 == opcode | 8'hf8 == opcode | 8'h58
     == opcode | 8'h78 == opcode | 8'hb8 == opcode | 8'hea == opcode ? regs_x : _GEN_1394; // @[CPU6502Core.scala 89:20 92:16]
  wire [7:0] execResult_result_1_regs_y = 8'h18 == opcode | 8'h38 == opcode | 8'hd8 == opcode | 8'hf8 == opcode | 8'h58
     == opcode | 8'h78 == opcode | 8'hb8 == opcode | 8'hea == opcode ? regs_y : _GEN_1395; // @[CPU6502Core.scala 89:20 92:16]
  wire [7:0] execResult_result_1_regs_sp = 8'h18 == opcode | 8'h38 == opcode | 8'hd8 == opcode | 8'hf8 == opcode | 8'h58
     == opcode | 8'h78 == opcode | 8'hb8 == opcode | 8'hea == opcode ? regs_sp : _GEN_1396; // @[CPU6502Core.scala 89:20 92:16]
  wire [15:0] execResult_result_1_regs_pc = 8'h18 == opcode | 8'h38 == opcode | 8'hd8 == opcode | 8'hf8 == opcode | 8'h58
     == opcode | 8'h78 == opcode | 8'hb8 == opcode | 8'hea == opcode ? regs_pc : _GEN_1397; // @[CPU6502Core.scala 89:20 92:16]
  wire  execResult_result_1_regs_flagC = 8'h18 == opcode | 8'h38 == opcode | 8'hd8 == opcode | 8'hf8 == opcode | 8'h58
     == opcode | 8'h78 == opcode | 8'hb8 == opcode | 8'hea == opcode ? execResult_result_newRegs_flagC : _GEN_1398; // @[CPU6502Core.scala 89:20 92:16]
  wire  execResult_result_1_regs_flagZ = 8'h18 == opcode | 8'h38 == opcode | 8'hd8 == opcode | 8'hf8 == opcode | 8'h58
     == opcode | 8'h78 == opcode | 8'hb8 == opcode | 8'hea == opcode ? regs_flagZ : _GEN_1399; // @[CPU6502Core.scala 89:20 92:16]
  wire  execResult_result_1_regs_flagI = 8'h18 == opcode | 8'h38 == opcode | 8'hd8 == opcode | 8'hf8 == opcode | 8'h58
     == opcode | 8'h78 == opcode | 8'hb8 == opcode | 8'hea == opcode ? execResult_result_newRegs_flagI : _GEN_1400; // @[CPU6502Core.scala 89:20 92:16]
  wire  execResult_result_1_regs_flagD = 8'h18 == opcode | 8'h38 == opcode | 8'hd8 == opcode | 8'hf8 == opcode | 8'h58
     == opcode | 8'h78 == opcode | 8'hb8 == opcode | 8'hea == opcode ? execResult_result_newRegs_flagD : _GEN_1401; // @[CPU6502Core.scala 89:20 92:16]
  wire  execResult_result_1_regs_flagV = 8'h18 == opcode | 8'h38 == opcode | 8'hd8 == opcode | 8'hf8 == opcode | 8'h58
     == opcode | 8'h78 == opcode | 8'hb8 == opcode | 8'hea == opcode ? execResult_result_newRegs_flagV : _GEN_1403; // @[CPU6502Core.scala 89:20 92:16]
  wire  execResult_result_1_regs_flagN = 8'h18 == opcode | 8'h38 == opcode | 8'hd8 == opcode | 8'hf8 == opcode | 8'h58
     == opcode | 8'h78 == opcode | 8'hb8 == opcode | 8'hea == opcode ? regs_flagN : _GEN_1404; // @[CPU6502Core.scala 89:20 92:16]
  wire [15:0] execResult_result_1_memAddr = 8'h18 == opcode | 8'h38 == opcode | 8'hd8 == opcode | 8'hf8 == opcode | 8'h58
     == opcode | 8'h78 == opcode | 8'hb8 == opcode | 8'hea == opcode ? 16'h0 : _GEN_1405; // @[CPU6502Core.scala 89:20 92:16]
  wire [7:0] execResult_result_1_memData = 8'h18 == opcode | 8'h38 == opcode | 8'hd8 == opcode | 8'hf8 == opcode | 8'h58
     == opcode | 8'h78 == opcode | 8'hb8 == opcode | 8'hea == opcode ? 8'h0 : _GEN_1406; // @[CPU6502Core.scala 89:20 92:16]
  wire  execResult_result_1_memWrite = 8'h18 == opcode | 8'h38 == opcode | 8'hd8 == opcode | 8'hf8 == opcode | 8'h58 ==
    opcode | 8'h78 == opcode | 8'hb8 == opcode | 8'hea == opcode ? 1'h0 : _GEN_1407; // @[CPU6502Core.scala 89:20 92:16]
  wire  execResult_result_1_memRead = 8'h18 == opcode | 8'h38 == opcode | 8'hd8 == opcode | 8'hf8 == opcode | 8'h58 ==
    opcode | 8'h78 == opcode | 8'hb8 == opcode | 8'hea == opcode ? 1'h0 : _GEN_1408; // @[CPU6502Core.scala 89:20 92:16]
  wire [15:0] execResult_result_1_operand = 8'h18 == opcode | 8'h38 == opcode | 8'hd8 == opcode | 8'hf8 == opcode | 8'h58
     == opcode | 8'h78 == opcode | 8'hb8 == opcode | 8'hea == opcode ? 16'h0 : _GEN_1409; // @[CPU6502Core.scala 89:20 92:16]
  wire  _GEN_1431 = 2'h1 == state & execResult_result_1_done; // @[CPU6502Core.scala 37:14 40:17 52:18]
  wire  execResult_done = 2'h0 == state ? 1'h0 : _GEN_1431; // @[CPU6502Core.scala 37:14 40:17]
  wire [2:0] _GEN_1432 = 2'h1 == state ? execResult_result_1_nextCycle : 3'h0; // @[CPU6502Core.scala 37:14 40:17 52:18]
  wire [2:0] execResult_nextCycle = 2'h0 == state ? 3'h0 : _GEN_1432; // @[CPU6502Core.scala 37:14 40:17]
  wire [7:0] _GEN_1433 = 2'h1 == state ? execResult_result_1_regs_a : regs_a; // @[CPU6502Core.scala 37:14 40:17 52:18]
  wire [7:0] _GEN_1434 = 2'h1 == state ? execResult_result_1_regs_x : regs_x; // @[CPU6502Core.scala 37:14 40:17 52:18]
  wire [7:0] _GEN_1435 = 2'h1 == state ? execResult_result_1_regs_y : regs_y; // @[CPU6502Core.scala 37:14 40:17 52:18]
  wire [7:0] _GEN_1436 = 2'h1 == state ? execResult_result_1_regs_sp : regs_sp; // @[CPU6502Core.scala 37:14 40:17 52:18]
  wire [15:0] _GEN_1437 = 2'h1 == state ? execResult_result_1_regs_pc : regs_pc; // @[CPU6502Core.scala 37:14 40:17 52:18]
  wire  _GEN_1438 = 2'h1 == state ? execResult_result_1_regs_flagC : regs_flagC; // @[CPU6502Core.scala 37:14 40:17 52:18]
  wire  _GEN_1439 = 2'h1 == state ? execResult_result_1_regs_flagZ : regs_flagZ; // @[CPU6502Core.scala 37:14 40:17 52:18]
  wire  _GEN_1440 = 2'h1 == state ? execResult_result_1_regs_flagI : regs_flagI; // @[CPU6502Core.scala 37:14 40:17 52:18]
  wire  _GEN_1441 = 2'h1 == state ? execResult_result_1_regs_flagD : regs_flagD; // @[CPU6502Core.scala 37:14 40:17 52:18]
  wire  _GEN_1443 = 2'h1 == state ? execResult_result_1_regs_flagV : regs_flagV; // @[CPU6502Core.scala 37:14 40:17 52:18]
  wire  _GEN_1444 = 2'h1 == state ? execResult_result_1_regs_flagN : regs_flagN; // @[CPU6502Core.scala 37:14 40:17 52:18]
  wire [15:0] _GEN_1445 = 2'h1 == state ? execResult_result_1_memAddr : 16'h0; // @[CPU6502Core.scala 37:14 40:17 52:18]
  wire [7:0] _GEN_1446 = 2'h1 == state ? execResult_result_1_memData : 8'h0; // @[CPU6502Core.scala 37:14 40:17 52:18]
  wire  _GEN_1447 = 2'h1 == state & execResult_result_1_memWrite; // @[CPU6502Core.scala 37:14 40:17 52:18]
  wire  _GEN_1448 = 2'h1 == state & execResult_result_1_memRead; // @[CPU6502Core.scala 37:14 40:17 52:18]
  wire [15:0] _GEN_1449 = 2'h1 == state ? execResult_result_1_operand : operand; // @[CPU6502Core.scala 37:14 40:17 52:18]
  wire [15:0] execResult_memAddr = 2'h0 == state ? 16'h0 : _GEN_1445; // @[CPU6502Core.scala 37:14 40:17]
  wire [15:0] _GEN_1450 = 2'h1 == state ? execResult_memAddr : regs_pc; // @[CPU6502Core.scala 30:17 40:17 55:21]
  wire [7:0] execResult_memData = 2'h0 == state ? 8'h0 : _GEN_1446; // @[CPU6502Core.scala 37:14 40:17]
  wire [7:0] _GEN_1451 = 2'h1 == state ? execResult_memData : 8'h0; // @[CPU6502Core.scala 31:17 40:17 56:21]
  wire  execResult_memWrite = 2'h0 == state ? 1'h0 : _GEN_1447; // @[CPU6502Core.scala 37:14 40:17]
  wire  _GEN_1452 = 2'h1 == state & execResult_memWrite; // @[CPU6502Core.scala 32:17 40:17 57:21]
  wire  execResult_memRead = 2'h0 == state ? 1'h0 : _GEN_1448; // @[CPU6502Core.scala 37:14 40:17]
  wire  _GEN_1453 = 2'h1 == state & execResult_memRead; // @[CPU6502Core.scala 33:17 40:17 58:21]
  assign io_memAddr = 2'h0 == state ? regs_pc : _GEN_1450; // @[CPU6502Core.scala 40:17 42:18]
  assign io_memDataOut = 2'h0 == state ? 8'h0 : _GEN_1451; // @[CPU6502Core.scala 31:17 40:17]
  assign io_memWrite = 2'h0 == state ? 1'h0 : _GEN_1452; // @[CPU6502Core.scala 32:17 40:17]
  assign io_memRead = 2'h0 == state | _GEN_1453; // @[CPU6502Core.scala 40:17 43:18]
  assign io_debug_regA = regs_a; // @[DebugBundle.scala 21:21 22:16]
  assign io_debug_regX = regs_x; // @[DebugBundle.scala 21:21 23:16]
  assign io_debug_regY = regs_y; // @[DebugBundle.scala 21:21 24:16]
  assign io_debug_regPC = regs_pc; // @[DebugBundle.scala 21:21 25:17]
  assign io_debug_regSP = regs_sp; // @[DebugBundle.scala 21:21 26:17]
  assign io_debug_flagC = regs_flagC; // @[DebugBundle.scala 21:21 27:17]
  assign io_debug_flagZ = regs_flagZ; // @[DebugBundle.scala 21:21 28:17]
  assign io_debug_flagN = regs_flagN; // @[DebugBundle.scala 21:21 29:17]
  assign io_debug_flagV = regs_flagV; // @[DebugBundle.scala 21:21 30:17]
  assign io_debug_opcode = opcode; // @[DebugBundle.scala 21:21 31:18]
  always @(posedge clock) begin
    if (reset) begin // @[CPU6502Core.scala 19:21]
      regs_a <= 8'h0; // @[CPU6502Core.scala 19:21]
    end else if (!(2'h0 == state)) begin // @[CPU6502Core.scala 40:17]
      if (2'h1 == state) begin // @[CPU6502Core.scala 40:17]
        if (!(2'h0 == state)) begin // @[CPU6502Core.scala 40:17]
          regs_a <= _GEN_1433;
        end
      end
    end
    if (reset) begin // @[CPU6502Core.scala 19:21]
      regs_x <= 8'h0; // @[CPU6502Core.scala 19:21]
    end else if (!(2'h0 == state)) begin // @[CPU6502Core.scala 40:17]
      if (2'h1 == state) begin // @[CPU6502Core.scala 40:17]
        if (!(2'h0 == state)) begin // @[CPU6502Core.scala 40:17]
          regs_x <= _GEN_1434;
        end
      end
    end
    if (reset) begin // @[CPU6502Core.scala 19:21]
      regs_y <= 8'h0; // @[CPU6502Core.scala 19:21]
    end else if (!(2'h0 == state)) begin // @[CPU6502Core.scala 40:17]
      if (2'h1 == state) begin // @[CPU6502Core.scala 40:17]
        if (!(2'h0 == state)) begin // @[CPU6502Core.scala 40:17]
          regs_y <= _GEN_1435;
        end
      end
    end
    if (reset) begin // @[CPU6502Core.scala 19:21]
      regs_sp <= 8'hff; // @[CPU6502Core.scala 19:21]
    end else if (!(2'h0 == state)) begin // @[CPU6502Core.scala 40:17]
      if (2'h1 == state) begin // @[CPU6502Core.scala 40:17]
        if (!(2'h0 == state)) begin // @[CPU6502Core.scala 40:17]
          regs_sp <= _GEN_1436;
        end
      end
    end
    if (reset) begin // @[CPU6502Core.scala 19:21]
      regs_pc <= 16'h0; // @[CPU6502Core.scala 19:21]
    end else if (2'h0 == state) begin // @[CPU6502Core.scala 40:17]
      regs_pc <= _regs_pc_T_1; // @[CPU6502Core.scala 45:15]
    end else if (2'h1 == state) begin // @[CPU6502Core.scala 40:17]
      if (!(2'h0 == state)) begin // @[CPU6502Core.scala 40:17]
        regs_pc <= _GEN_1437;
      end
    end
    if (reset) begin // @[CPU6502Core.scala 19:21]
      regs_flagC <= 1'h0; // @[CPU6502Core.scala 19:21]
    end else if (!(2'h0 == state)) begin // @[CPU6502Core.scala 40:17]
      if (2'h1 == state) begin // @[CPU6502Core.scala 40:17]
        if (!(2'h0 == state)) begin // @[CPU6502Core.scala 40:17]
          regs_flagC <= _GEN_1438;
        end
      end
    end
    if (reset) begin // @[CPU6502Core.scala 19:21]
      regs_flagZ <= 1'h0; // @[CPU6502Core.scala 19:21]
    end else if (!(2'h0 == state)) begin // @[CPU6502Core.scala 40:17]
      if (2'h1 == state) begin // @[CPU6502Core.scala 40:17]
        if (!(2'h0 == state)) begin // @[CPU6502Core.scala 40:17]
          regs_flagZ <= _GEN_1439;
        end
      end
    end
    if (reset) begin // @[CPU6502Core.scala 19:21]
      regs_flagI <= 1'h0; // @[CPU6502Core.scala 19:21]
    end else if (!(2'h0 == state)) begin // @[CPU6502Core.scala 40:17]
      if (2'h1 == state) begin // @[CPU6502Core.scala 40:17]
        if (!(2'h0 == state)) begin // @[CPU6502Core.scala 40:17]
          regs_flagI <= _GEN_1440;
        end
      end
    end
    if (reset) begin // @[CPU6502Core.scala 19:21]
      regs_flagD <= 1'h0; // @[CPU6502Core.scala 19:21]
    end else if (!(2'h0 == state)) begin // @[CPU6502Core.scala 40:17]
      if (2'h1 == state) begin // @[CPU6502Core.scala 40:17]
        if (!(2'h0 == state)) begin // @[CPU6502Core.scala 40:17]
          regs_flagD <= _GEN_1441;
        end
      end
    end
    if (reset) begin // @[CPU6502Core.scala 19:21]
      regs_flagV <= 1'h0; // @[CPU6502Core.scala 19:21]
    end else if (!(2'h0 == state)) begin // @[CPU6502Core.scala 40:17]
      if (2'h1 == state) begin // @[CPU6502Core.scala 40:17]
        if (!(2'h0 == state)) begin // @[CPU6502Core.scala 40:17]
          regs_flagV <= _GEN_1443;
        end
      end
    end
    if (reset) begin // @[CPU6502Core.scala 19:21]
      regs_flagN <= 1'h0; // @[CPU6502Core.scala 19:21]
    end else if (!(2'h0 == state)) begin // @[CPU6502Core.scala 40:17]
      if (2'h1 == state) begin // @[CPU6502Core.scala 40:17]
        if (!(2'h0 == state)) begin // @[CPU6502Core.scala 40:17]
          regs_flagN <= _GEN_1444;
        end
      end
    end
    if (reset) begin // @[CPU6502Core.scala 23:22]
      state <= 2'h0; // @[CPU6502Core.scala 23:22]
    end else if (2'h0 == state) begin // @[CPU6502Core.scala 40:17]
      state <= 2'h1; // @[CPU6502Core.scala 47:13]
    end else if (2'h1 == state) begin // @[CPU6502Core.scala 40:17]
      if (execResult_done) begin // @[CPU6502Core.scala 64:29]
        state <= 2'h0; // @[CPU6502Core.scala 66:15]
      end
    end
    if (reset) begin // @[CPU6502Core.scala 25:24]
      opcode <= 8'h0; // @[CPU6502Core.scala 25:24]
    end else if (2'h0 == state) begin // @[CPU6502Core.scala 40:17]
      opcode <= io_memDataIn; // @[CPU6502Core.scala 44:14]
    end
    if (reset) begin // @[CPU6502Core.scala 26:24]
      operand <= 16'h0; // @[CPU6502Core.scala 26:24]
    end else if (!(2'h0 == state)) begin // @[CPU6502Core.scala 40:17]
      if (2'h1 == state) begin // @[CPU6502Core.scala 40:17]
        if (!(2'h0 == state)) begin // @[CPU6502Core.scala 40:17]
          operand <= _GEN_1449;
        end
      end
    end
    if (reset) begin // @[CPU6502Core.scala 27:24]
      cycle <= 3'h0; // @[CPU6502Core.scala 27:24]
    end else if (2'h0 == state) begin // @[CPU6502Core.scala 40:17]
      cycle <= 3'h0; // @[CPU6502Core.scala 46:13]
    end else if (2'h1 == state) begin // @[CPU6502Core.scala 40:17]
      if (execResult_done) begin // @[CPU6502Core.scala 64:29]
        cycle <= 3'h0; // @[CPU6502Core.scala 65:15]
      end else begin
        cycle <= execResult_nextCycle; // @[CPU6502Core.scala 62:15]
      end
    end
  end
endmodule
module CPU6502Refactored(
  input         clock,
  input         reset,
  output [15:0] io_memAddr,
  output [7:0]  io_memDataOut,
  input  [7:0]  io_memDataIn,
  output        io_memWrite,
  output        io_memRead,
  output [7:0]  io_debug_regA,
  output [7:0]  io_debug_regX,
  output [7:0]  io_debug_regY,
  output [15:0] io_debug_regPC,
  output [7:0]  io_debug_regSP,
  output        io_debug_flagC,
  output        io_debug_flagZ,
  output        io_debug_flagN,
  output        io_debug_flagV,
  output [7:0]  io_debug_opcode
);
  wire  core_clock; // @[CPU6502Refactored.scala 18:20]
  wire  core_reset; // @[CPU6502Refactored.scala 18:20]
  wire [15:0] core_io_memAddr; // @[CPU6502Refactored.scala 18:20]
  wire [7:0] core_io_memDataOut; // @[CPU6502Refactored.scala 18:20]
  wire [7:0] core_io_memDataIn; // @[CPU6502Refactored.scala 18:20]
  wire  core_io_memWrite; // @[CPU6502Refactored.scala 18:20]
  wire  core_io_memRead; // @[CPU6502Refactored.scala 18:20]
  wire [7:0] core_io_debug_regA; // @[CPU6502Refactored.scala 18:20]
  wire [7:0] core_io_debug_regX; // @[CPU6502Refactored.scala 18:20]
  wire [7:0] core_io_debug_regY; // @[CPU6502Refactored.scala 18:20]
  wire [15:0] core_io_debug_regPC; // @[CPU6502Refactored.scala 18:20]
  wire [7:0] core_io_debug_regSP; // @[CPU6502Refactored.scala 18:20]
  wire  core_io_debug_flagC; // @[CPU6502Refactored.scala 18:20]
  wire  core_io_debug_flagZ; // @[CPU6502Refactored.scala 18:20]
  wire  core_io_debug_flagN; // @[CPU6502Refactored.scala 18:20]
  wire  core_io_debug_flagV; // @[CPU6502Refactored.scala 18:20]
  wire [7:0] core_io_debug_opcode; // @[CPU6502Refactored.scala 18:20]
  CPU6502Core core ( // @[CPU6502Refactored.scala 18:20]
    .clock(core_clock),
    .reset(core_reset),
    .io_memAddr(core_io_memAddr),
    .io_memDataOut(core_io_memDataOut),
    .io_memDataIn(core_io_memDataIn),
    .io_memWrite(core_io_memWrite),
    .io_memRead(core_io_memRead),
    .io_debug_regA(core_io_debug_regA),
    .io_debug_regX(core_io_debug_regX),
    .io_debug_regY(core_io_debug_regY),
    .io_debug_regPC(core_io_debug_regPC),
    .io_debug_regSP(core_io_debug_regSP),
    .io_debug_flagC(core_io_debug_flagC),
    .io_debug_flagZ(core_io_debug_flagZ),
    .io_debug_flagN(core_io_debug_flagN),
    .io_debug_flagV(core_io_debug_flagV),
    .io_debug_opcode(core_io_debug_opcode)
  );
  assign io_memAddr = core_io_memAddr; // @[CPU6502Refactored.scala 20:17]
  assign io_memDataOut = core_io_memDataOut; // @[CPU6502Refactored.scala 21:17]
  assign io_memWrite = core_io_memWrite; // @[CPU6502Refactored.scala 23:17]
  assign io_memRead = core_io_memRead; // @[CPU6502Refactored.scala 24:17]
  assign io_debug_regA = core_io_debug_regA; // @[CPU6502Refactored.scala 25:17]
  assign io_debug_regX = core_io_debug_regX; // @[CPU6502Refactored.scala 25:17]
  assign io_debug_regY = core_io_debug_regY; // @[CPU6502Refactored.scala 25:17]
  assign io_debug_regPC = core_io_debug_regPC; // @[CPU6502Refactored.scala 25:17]
  assign io_debug_regSP = core_io_debug_regSP; // @[CPU6502Refactored.scala 25:17]
  assign io_debug_flagC = core_io_debug_flagC; // @[CPU6502Refactored.scala 25:17]
  assign io_debug_flagZ = core_io_debug_flagZ; // @[CPU6502Refactored.scala 25:17]
  assign io_debug_flagN = core_io_debug_flagN; // @[CPU6502Refactored.scala 25:17]
  assign io_debug_flagV = core_io_debug_flagV; // @[CPU6502Refactored.scala 25:17]
  assign io_debug_opcode = core_io_debug_opcode; // @[CPU6502Refactored.scala 25:17]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_memDataIn = io_memDataIn; // @[CPU6502Refactored.scala 22:21]
endmodule
