module CPU6502(
  input         clock,
  input         reset,
  output [15:0] io_memAddr,
  output [7:0]  io_memDataOut,
  input  [7:0]  io_memDataIn,
  output        io_memWrite,
  output        io_memRead,
  output [7:0]  io_debug_regA,
  output [7:0]  io_debug_regX,
  output [7:0]  io_debug_regY,
  output [15:0] io_debug_regPC,
  output [7:0]  io_debug_regSP,
  output        io_debug_flagC,
  output        io_debug_flagZ,
  output        io_debug_flagN,
  output        io_debug_flagV,
  output [7:0]  io_debug_opcode
);
  reg [7:0] regA; // @[CPU6502.scala 18:21]
  reg [7:0] regX; // @[CPU6502.scala 19:21]
  reg [7:0] regY; // @[CPU6502.scala 20:21]
  reg [7:0] regSP; // @[CPU6502.scala 21:22]
  reg [15:0] regPC; // @[CPU6502.scala 22:22]
  reg  flagC; // @[CPU6502.scala 25:22]
  reg  flagZ; // @[CPU6502.scala 26:22]
  reg  flagI; // @[CPU6502.scala 27:22]
  reg  flagD; // @[CPU6502.scala 28:22]
  reg  flagV; // @[CPU6502.scala 30:22]
  reg  flagN; // @[CPU6502.scala 31:22]
  reg [1:0] state; // @[CPU6502.scala 35:22]
  reg [7:0] opcode; // @[CPU6502.scala 37:23]
  reg [15:0] operand; // @[CPU6502.scala 38:24]
  reg [2:0] cycle; // @[CPU6502.scala 39:22]
  wire [15:0] _regPC_T_1 = regPC + 16'h1; // @[CPU6502.scala 60:22]
  wire  _T_3 = cycle == 3'h0; // @[CPU6502.scala 69:22]
  wire [7:0] _GEN_2 = cycle == 3'h0 ? io_memDataIn : regA; // @[CPU6502.scala 69:31 72:18 18:21]
  wire  _GEN_3 = cycle == 3'h0 ? io_memDataIn[7] : flagN; // @[CPU6502.scala 50:11 31:22 69:31]
  wire  _GEN_4 = cycle == 3'h0 ? io_memDataIn == 8'h0 : flagZ; // @[CPU6502.scala 51:11 26:22 69:31]
  wire [15:0] _GEN_5 = cycle == 3'h0 ? _regPC_T_1 : regPC; // @[CPU6502.scala 69:31 74:19 22:22]
  wire [1:0] _GEN_6 = cycle == 3'h0 ? 2'h0 : state; // @[CPU6502.scala 69:31 75:19 35:22]
  wire  _T_6 = cycle == 3'h1; // @[CPU6502.scala 86:28]
  wire [15:0] _GEN_7 = cycle == 3'h1 ? operand : regPC; // @[CPU6502.scala 42:14 86:37 87:24]
  wire [7:0] _GEN_9 = cycle == 3'h1 ? io_memDataIn : regA; // @[CPU6502.scala 86:37 89:18 18:21]
  wire  _GEN_10 = cycle == 3'h1 ? io_memDataIn[7] : flagN; // @[CPU6502.scala 50:11 31:22 86:37]
  wire  _GEN_11 = cycle == 3'h1 ? io_memDataIn == 8'h0 : flagZ; // @[CPU6502.scala 51:11 26:22 86:37]
  wire [1:0] _GEN_12 = cycle == 3'h1 ? 2'h0 : state; // @[CPU6502.scala 86:37 91:19 35:22]
  wire [15:0] _GEN_13 = _T_3 ? regPC : _GEN_7; // @[CPU6502.scala 80:31 81:24]
  wire  _GEN_14 = _T_3 | _T_6; // @[CPU6502.scala 80:31 82:24]
  wire [15:0] _GEN_15 = _T_3 ? {{8'd0}, io_memDataIn} : operand; // @[CPU6502.scala 80:31 83:21 38:24]
  wire [2:0] _GEN_17 = _T_3 ? 3'h1 : cycle; // @[CPU6502.scala 80:31 85:19 39:22]
  wire [7:0] _GEN_18 = _T_3 ? regA : _GEN_9; // @[CPU6502.scala 18:21 80:31]
  wire  _GEN_19 = _T_3 ? flagN : _GEN_10; // @[CPU6502.scala 31:22 80:31]
  wire  _GEN_20 = _T_3 ? flagZ : _GEN_11; // @[CPU6502.scala 26:22 80:31]
  wire [1:0] _GEN_21 = _T_3 ? state : _GEN_12; // @[CPU6502.scala 35:22 80:31]
  wire [7:0] _GEN_24 = _T_3 ? io_memDataIn : regX; // @[CPU6502.scala 100:18 19:21 97:31]
  wire [7:0] _GEN_31 = _T_3 ? io_memDataIn : regY; // @[CPU6502.scala 109:31 112:18 20:21]
  wire [7:0] _GEN_37 = _T_6 ? regA : 8'h0; // @[CPU6502.scala 127:37 129:27 43:17]
  wire [7:0] _GEN_45 = _T_3 ? 8'h0 : _GEN_37; // @[CPU6502.scala 121:31 43:17]
  wire  _GEN_46 = _T_3 ? 1'h0 : _T_6; // @[CPU6502.scala 121:31 44:15]
  wire [8:0] _sum_T = regA + io_memDataIn; // @[CPU6502.scala 140:28]
  wire [8:0] _GEN_1892 = {{8'd0}, flagC}; // @[CPU6502.scala 140:44]
  wire [9:0] sum = _sum_T + _GEN_1892; // @[CPU6502.scala 140:44]
  wire [7:0] sum8 = sum[7:0]; // @[CPU6502.scala 141:27]
  wire [7:0] _GEN_50 = _T_3 ? sum8 : regA; // @[CPU6502.scala 137:31 142:18 18:21]
  wire  _GEN_51 = _T_3 ? sum[8] : flagC; // @[CPU6502.scala 137:31 143:19 25:22]
  wire  _GEN_52 = _T_3 ? sum8[7] : flagN; // @[CPU6502.scala 137:31 50:11 31:22]
  wire  _GEN_53 = _T_3 ? sum8 == 8'h0 : flagZ; // @[CPU6502.scala 137:31 51:11 26:22]
  wire  _GEN_54 = _T_3 ? regA[7] == io_memDataIn[7] & regA[7] != sum[7] : flagV; // @[CPU6502.scala 137:31 146:19 30:22]
  wire [8:0] _diff_T = regA - io_memDataIn; // @[CPU6502.scala 157:29]
  wire  _diff_T_2 = ~flagC; // @[CPU6502.scala 157:49]
  wire [8:0] _GEN_1893 = {{8'd0}, _diff_T_2}; // @[CPU6502.scala 157:45]
  wire [9:0] diff = _diff_T - _GEN_1893; // @[CPU6502.scala 157:45]
  wire [7:0] diff8 = diff[7:0]; // @[CPU6502.scala 158:29]
  wire [7:0] _GEN_59 = _T_3 ? diff8 : regA; // @[CPU6502.scala 154:31 159:18 18:21]
  wire  _GEN_60 = _T_3 ? ~diff[8] : flagC; // @[CPU6502.scala 154:31 160:19 25:22]
  wire  _GEN_61 = _T_3 ? diff8[7] : flagN; // @[CPU6502.scala 154:31 50:11 31:22]
  wire  _GEN_62 = _T_3 ? diff8 == 8'h0 : flagZ; // @[CPU6502.scala 154:31 51:11 26:22]
  wire  _GEN_63 = _T_3 ? regA[7] != io_memDataIn[7] & regA[7] != diff[7] : flagV; // @[CPU6502.scala 154:31 162:19 30:22]
  wire [7:0] result = regA & io_memDataIn; // @[CPU6502.scala 173:31]
  wire  _flagZ_T_6 = result == 8'h0; // @[CPU6502.scala 51:20]
  wire [7:0] _GEN_68 = _T_3 ? result : regA; // @[CPU6502.scala 170:31 174:18 18:21]
  wire  _GEN_69 = _T_3 ? result[7] : flagN; // @[CPU6502.scala 170:31 50:11 31:22]
  wire  _GEN_70 = _T_3 ? result == 8'h0 : flagZ; // @[CPU6502.scala 170:31 51:11 26:22]
  wire [7:0] result_1 = regA | io_memDataIn; // @[CPU6502.scala 186:31]
  wire [7:0] _GEN_75 = _T_3 ? result_1 : regA; // @[CPU6502.scala 183:31 187:18 18:21]
  wire  _GEN_76 = _T_3 ? result_1[7] : flagN; // @[CPU6502.scala 183:31 50:11 31:22]
  wire  _GEN_77 = _T_3 ? result_1 == 8'h0 : flagZ; // @[CPU6502.scala 183:31 51:11 26:22]
  wire [7:0] result_2 = regA ^ io_memDataIn; // @[CPU6502.scala 199:31]
  wire [7:0] _GEN_82 = _T_3 ? result_2 : regA; // @[CPU6502.scala 196:31 200:18 18:21]
  wire  _GEN_83 = _T_3 ? result_2[7] : flagN; // @[CPU6502.scala 196:31 50:11 31:22]
  wire  _GEN_84 = _T_3 ? result_2 == 8'h0 : flagZ; // @[CPU6502.scala 196:31 51:11 26:22]
  wire [7:0] result_3 = regX + 8'h1; // @[CPU6502.scala 209:29]
  wire [7:0] result_4 = regY + 8'h1; // @[CPU6502.scala 217:29]
  wire [7:0] result_5 = regX - 8'h1; // @[CPU6502.scala 225:29]
  wire [7:0] result_6 = regY - 8'h1; // @[CPU6502.scala 233:29]
  wire [15:0] _regPC_T_25 = {io_memDataIn,operand[7:0]}; // @[Cat.scala 33:92]
  wire [15:0] _GEN_89 = _T_6 ? _regPC_T_25 : regPC; // @[CPU6502.scala 322:37 325:19 22:22]
  wire [15:0] _GEN_94 = _T_3 ? _regPC_T_1 : _GEN_89; // @[CPU6502.scala 316:31 320:19]
  wire [7:0] offset = io_memDataIn; // @[CPU6502.scala 337:41]
  wire [15:0] _GEN_1894 = {{8{offset[7]}},offset}; // @[CPU6502.scala 338:38]
  wire [15:0] _regPC_T_32 = $signed(regPC) + $signed(_GEN_1894); // @[CPU6502.scala 338:48]
  wire [15:0] _GEN_97 = flagZ ? _regPC_T_32 : _regPC_T_1; // @[CPU6502.scala 335:19 336:25 338:21]
  wire [15:0] _GEN_100 = _T_3 ? _GEN_97 : regPC; // @[CPU6502.scala 22:22 332:31]
  wire [15:0] _GEN_102 = ~flagZ ? _regPC_T_32 : _regPC_T_1; // @[CPU6502.scala 349:19 350:26 352:21]
  wire [15:0] _GEN_105 = _T_3 ? _GEN_102 : regPC; // @[CPU6502.scala 22:22 346:31]
  wire [15:0] _GEN_107 = flagC ? _regPC_T_32 : _regPC_T_1; // @[CPU6502.scala 363:19 364:25 366:21]
  wire [15:0] _GEN_110 = _T_3 ? _GEN_107 : regPC; // @[CPU6502.scala 22:22 360:31]
  wire [15:0] _GEN_112 = _diff_T_2 ? _regPC_T_32 : _regPC_T_1; // @[CPU6502.scala 377:19 378:26 380:21]
  wire [15:0] _GEN_115 = _T_3 ? _GEN_112 : regPC; // @[CPU6502.scala 22:22 374:31]
  wire [15:0] _GEN_117 = flagN ? _regPC_T_32 : _regPC_T_1; // @[CPU6502.scala 391:19 392:25 394:21]
  wire [15:0] _GEN_120 = _T_3 ? _GEN_117 : regPC; // @[CPU6502.scala 22:22 388:31]
  wire [15:0] _GEN_122 = ~flagN ? _regPC_T_32 : _regPC_T_1; // @[CPU6502.scala 405:19 406:26 408:21]
  wire [15:0] _GEN_125 = _T_3 ? _GEN_122 : regPC; // @[CPU6502.scala 22:22 402:31]
  wire [15:0] _GEN_127 = ~flagV ? _regPC_T_32 : _regPC_T_1; // @[CPU6502.scala 419:19 420:26 422:21]
  wire [15:0] _GEN_130 = _T_3 ? _GEN_127 : regPC; // @[CPU6502.scala 22:22 416:31]
  wire [15:0] _GEN_132 = flagV ? _regPC_T_32 : _regPC_T_1; // @[CPU6502.scala 433:19 434:25 436:21]
  wire [15:0] _GEN_135 = _T_3 ? _GEN_132 : regPC; // @[CPU6502.scala 22:22 430:31]
  wire  _flagC_T_3 = regA >= io_memDataIn; // @[CPU6502.scala 448:27]
  wire  _flagZ_T_17 = regA == io_memDataIn; // @[CPU6502.scala 449:27]
  wire  _GEN_139 = _T_3 ? regA >= io_memDataIn : flagC; // @[CPU6502.scala 444:31 448:19 25:22]
  wire  _GEN_140 = _T_3 ? regA == io_memDataIn : flagZ; // @[CPU6502.scala 444:31 449:19 26:22]
  wire  _GEN_141 = _T_3 ? _diff_T[7] : flagN; // @[CPU6502.scala 444:31 450:19 31:22]
  wire  _GEN_146 = _T_6 ? _flagC_T_3 : flagC; // @[CPU6502.scala 464:37 468:19 25:22]
  wire  _GEN_147 = _T_6 ? _flagZ_T_17 : flagZ; // @[CPU6502.scala 464:37 469:19 26:22]
  wire  _GEN_148 = _T_6 ? _diff_T[7] : flagN; // @[CPU6502.scala 464:37 470:19 31:22]
  wire  _GEN_155 = _T_3 ? flagC : _GEN_146; // @[CPU6502.scala 25:22 458:31]
  wire  _GEN_156 = _T_3 ? flagZ : _GEN_147; // @[CPU6502.scala 26:22 458:31]
  wire  _GEN_157 = _T_3 ? flagN : _GEN_148; // @[CPU6502.scala 31:22 458:31]
  wire [8:0] result_9 = regX - io_memDataIn; // @[CPU6502.scala 480:31]
  wire  _GEN_161 = _T_3 ? regX >= io_memDataIn : flagC; // @[CPU6502.scala 477:31 481:19 25:22]
  wire  _GEN_162 = _T_3 ? regX == io_memDataIn : flagZ; // @[CPU6502.scala 477:31 482:19 26:22]
  wire  _GEN_163 = _T_3 ? result_9[7] : flagN; // @[CPU6502.scala 477:31 483:19 31:22]
  wire [8:0] result_10 = regY - io_memDataIn; // @[CPU6502.scala 494:31]
  wire  _GEN_168 = _T_3 ? regY >= io_memDataIn : flagC; // @[CPU6502.scala 491:31 495:19 25:22]
  wire  _GEN_169 = _T_3 ? regY == io_memDataIn : flagZ; // @[CPU6502.scala 491:31 496:19 26:22]
  wire  _GEN_170 = _T_3 ? result_10[7] : flagN; // @[CPU6502.scala 491:31 497:19 31:22]
  wire  _GEN_175 = _T_6 ? _flagZ_T_6 : flagZ; // @[CPU6502.scala 511:37 515:19 26:22]
  wire  _GEN_177 = _T_6 ? io_memDataIn[6] : flagV; // @[CPU6502.scala 511:37 517:19 30:22]
  wire  _GEN_184 = _T_3 ? flagZ : _GEN_175; // @[CPU6502.scala 26:22 505:31]
  wire  _GEN_186 = _T_3 ? flagV : _GEN_177; // @[CPU6502.scala 30:22 505:31]
  wire [8:0] _result_T_8 = {regA, 1'h0}; // @[CPU6502.scala 526:27]
  wire [7:0] result_11 = _result_T_8[7:0]; // @[CPU6502.scala 526:32]
  wire  _T_79 = cycle == 3'h2; // @[CPU6502.scala 544:28]
  wire [7:0] result_12 = {io_memDataIn[6:0],1'h0}; // @[Cat.scala 33:92]
  wire [15:0] _GEN_188 = cycle == 3'h2 ? operand : regPC; // @[CPU6502.scala 42:14 544:37 545:24]
  wire  _GEN_189 = cycle == 3'h2 ? io_memDataIn[7] : flagC; // @[CPU6502.scala 544:37 547:19 25:22]
  wire [7:0] _GEN_190 = cycle == 3'h2 ? result_12 : 8'h0; // @[CPU6502.scala 43:17 544:37 549:27]
  wire  _GEN_192 = cycle == 3'h2 ? result_12[7] : flagN; // @[CPU6502.scala 50:11 31:22 544:37]
  wire  _GEN_193 = cycle == 3'h2 ? result_12 == 8'h0 : flagZ; // @[CPU6502.scala 51:11 26:22 544:37]
  wire [1:0] _GEN_194 = cycle == 3'h2 ? 2'h0 : state; // @[CPU6502.scala 544:37 552:19 35:22]
  wire [15:0] _GEN_195 = _T_6 ? operand : _GEN_188; // @[CPU6502.scala 540:37 541:24]
  wire [2:0] _GEN_197 = _T_6 ? 3'h2 : cycle; // @[CPU6502.scala 540:37 543:19 39:22]
  wire  _GEN_198 = _T_6 ? flagC : _GEN_189; // @[CPU6502.scala 25:22 540:37]
  wire [7:0] _GEN_199 = _T_6 ? 8'h0 : _GEN_190; // @[CPU6502.scala 43:17 540:37]
  wire  _GEN_200 = _T_6 ? 1'h0 : _T_79; // @[CPU6502.scala 44:15 540:37]
  wire  _GEN_201 = _T_6 ? flagN : _GEN_192; // @[CPU6502.scala 31:22 540:37]
  wire  _GEN_202 = _T_6 ? flagZ : _GEN_193; // @[CPU6502.scala 26:22 540:37]
  wire [1:0] _GEN_203 = _T_6 ? state : _GEN_194; // @[CPU6502.scala 35:22 540:37]
  wire [15:0] _GEN_204 = _T_3 ? regPC : _GEN_195; // @[CPU6502.scala 534:31 535:24]
  wire [2:0] _GEN_208 = _T_3 ? 3'h1 : _GEN_197; // @[CPU6502.scala 534:31 539:19]
  wire  _GEN_209 = _T_3 ? flagC : _GEN_198; // @[CPU6502.scala 25:22 534:31]
  wire [7:0] _GEN_210 = _T_3 ? 8'h0 : _GEN_199; // @[CPU6502.scala 43:17 534:31]
  wire  _GEN_211 = _T_3 ? 1'h0 : _GEN_200; // @[CPU6502.scala 44:15 534:31]
  wire  _GEN_212 = _T_3 ? flagN : _GEN_201; // @[CPU6502.scala 31:22 534:31]
  wire  _GEN_213 = _T_3 ? flagZ : _GEN_202; // @[CPU6502.scala 26:22 534:31]
  wire [1:0] _GEN_214 = _T_3 ? state : _GEN_203; // @[CPU6502.scala 35:22 534:31]
  wire [7:0] result_13 = {1'h0,regA[7:1]}; // @[Cat.scala 33:92]
  wire [7:0] result_14 = {1'h0,io_memDataIn[7:1]}; // @[Cat.scala 33:92]
  wire  _GEN_216 = _T_79 ? io_memDataIn[0] : flagC; // @[CPU6502.scala 577:37 580:19 25:22]
  wire [7:0] _GEN_217 = _T_79 ? result_14 : 8'h0; // @[CPU6502.scala 43:17 577:37 582:27]
  wire  _GEN_219 = _T_79 ? result_14[7] : flagN; // @[CPU6502.scala 50:11 31:22 577:37]
  wire  _GEN_220 = _T_79 ? result_14 == 8'h0 : flagZ; // @[CPU6502.scala 51:11 26:22 577:37]
  wire  _GEN_225 = _T_6 ? flagC : _GEN_216; // @[CPU6502.scala 25:22 573:37]
  wire [7:0] _GEN_226 = _T_6 ? 8'h0 : _GEN_217; // @[CPU6502.scala 43:17 573:37]
  wire  _GEN_228 = _T_6 ? flagN : _GEN_219; // @[CPU6502.scala 31:22 573:37]
  wire  _GEN_229 = _T_6 ? flagZ : _GEN_220; // @[CPU6502.scala 26:22 573:37]
  wire  _GEN_236 = _T_3 ? flagC : _GEN_225; // @[CPU6502.scala 25:22 567:31]
  wire [7:0] _GEN_237 = _T_3 ? 8'h0 : _GEN_226; // @[CPU6502.scala 43:17 567:31]
  wire  _GEN_239 = _T_3 ? flagN : _GEN_228; // @[CPU6502.scala 31:22 567:31]
  wire  _GEN_240 = _T_3 ? flagZ : _GEN_229; // @[CPU6502.scala 26:22 567:31]
  wire [7:0] result_15 = {regA[6:0],flagC}; // @[Cat.scala 33:92]
  wire [7:0] result_16 = {io_memDataIn[6:0],flagC}; // @[Cat.scala 33:92]
  wire [7:0] _GEN_244 = _T_79 ? result_16 : 8'h0; // @[CPU6502.scala 43:17 611:37 617:27]
  wire  _GEN_246 = _T_79 ? result_16[7] : flagN; // @[CPU6502.scala 50:11 31:22 611:37]
  wire  _GEN_247 = _T_79 ? result_16 == 8'h0 : flagZ; // @[CPU6502.scala 51:11 26:22 611:37]
  wire [7:0] _GEN_253 = _T_6 ? 8'h0 : _GEN_244; // @[CPU6502.scala 43:17 607:37]
  wire  _GEN_255 = _T_6 ? flagN : _GEN_246; // @[CPU6502.scala 31:22 607:37]
  wire  _GEN_256 = _T_6 ? flagZ : _GEN_247; // @[CPU6502.scala 26:22 607:37]
  wire [7:0] _GEN_264 = _T_3 ? 8'h0 : _GEN_253; // @[CPU6502.scala 43:17 601:31]
  wire  _GEN_266 = _T_3 ? flagN : _GEN_255; // @[CPU6502.scala 31:22 601:31]
  wire  _GEN_267 = _T_3 ? flagZ : _GEN_256; // @[CPU6502.scala 26:22 601:31]
  wire [7:0] result_17 = {flagC,regA[7:1]}; // @[Cat.scala 33:92]
  wire [7:0] result_18 = {flagC,io_memDataIn[7:1]}; // @[Cat.scala 33:92]
  wire [7:0] _GEN_271 = _T_79 ? result_18 : 8'h0; // @[CPU6502.scala 43:17 646:37 652:27]
  wire  _GEN_273 = _T_79 ? result_18[7] : flagN; // @[CPU6502.scala 50:11 31:22 646:37]
  wire  _GEN_274 = _T_79 ? result_18 == 8'h0 : flagZ; // @[CPU6502.scala 51:11 26:22 646:37]
  wire [7:0] _GEN_280 = _T_6 ? 8'h0 : _GEN_271; // @[CPU6502.scala 43:17 642:37]
  wire  _GEN_282 = _T_6 ? flagN : _GEN_273; // @[CPU6502.scala 31:22 642:37]
  wire  _GEN_283 = _T_6 ? flagZ : _GEN_274; // @[CPU6502.scala 26:22 642:37]
  wire [7:0] _GEN_291 = _T_3 ? 8'h0 : _GEN_280; // @[CPU6502.scala 43:17 636:31]
  wire  _GEN_293 = _T_3 ? flagN : _GEN_282; // @[CPU6502.scala 31:22 636:31]
  wire  _GEN_294 = _T_3 ? flagZ : _GEN_283; // @[CPU6502.scala 26:22 636:31]
  wire [7:0] result_19 = io_memDataIn + 8'h1; // @[CPU6502.scala 673:39]
  wire [7:0] _GEN_297 = _T_79 ? result_19 : 8'h0; // @[CPU6502.scala 43:17 671:37 674:27]
  wire  _GEN_299 = _T_79 ? result_19[7] : flagN; // @[CPU6502.scala 50:11 31:22 671:37]
  wire  _GEN_300 = _T_79 ? result_19 == 8'h0 : flagZ; // @[CPU6502.scala 51:11 26:22 671:37]
  wire [7:0] _GEN_305 = _T_6 ? 8'h0 : _GEN_297; // @[CPU6502.scala 43:17 667:37]
  wire  _GEN_307 = _T_6 ? flagN : _GEN_299; // @[CPU6502.scala 31:22 667:37]
  wire  _GEN_308 = _T_6 ? flagZ : _GEN_300; // @[CPU6502.scala 26:22 667:37]
  wire [7:0] _GEN_315 = _T_3 ? 8'h0 : _GEN_305; // @[CPU6502.scala 43:17 661:31]
  wire  _GEN_317 = _T_3 ? flagN : _GEN_307; // @[CPU6502.scala 31:22 661:31]
  wire  _GEN_318 = _T_3 ? flagZ : _GEN_308; // @[CPU6502.scala 26:22 661:31]
  wire [7:0] result_20 = io_memDataIn - 8'h1; // @[CPU6502.scala 695:39]
  wire [7:0] _GEN_321 = _T_79 ? result_20 : 8'h0; // @[CPU6502.scala 43:17 693:37 696:27]
  wire  _GEN_323 = _T_79 ? result_20[7] : flagN; // @[CPU6502.scala 50:11 31:22 693:37]
  wire  _GEN_324 = _T_79 ? result_20 == 8'h0 : flagZ; // @[CPU6502.scala 51:11 26:22 693:37]
  wire [7:0] _GEN_329 = _T_6 ? 8'h0 : _GEN_321; // @[CPU6502.scala 43:17 689:37]
  wire  _GEN_331 = _T_6 ? flagN : _GEN_323; // @[CPU6502.scala 31:22 689:37]
  wire  _GEN_332 = _T_6 ? flagZ : _GEN_324; // @[CPU6502.scala 26:22 689:37]
  wire [7:0] _GEN_339 = _T_3 ? 8'h0 : _GEN_329; // @[CPU6502.scala 43:17 683:31]
  wire  _GEN_341 = _T_3 ? flagN : _GEN_331; // @[CPU6502.scala 31:22 683:31]
  wire  _GEN_342 = _T_3 ? flagZ : _GEN_332; // @[CPU6502.scala 26:22 683:31]
  wire [7:0] _GEN_345 = _T_6 ? regX : 8'h0; // @[CPU6502.scala 43:17 711:37 713:27]
  wire [7:0] _GEN_353 = _T_3 ? 8'h0 : _GEN_345; // @[CPU6502.scala 43:17 705:31]
  wire [7:0] _GEN_357 = _T_6 ? regY : 8'h0; // @[CPU6502.scala 43:17 727:37 729:27]
  wire [7:0] _GEN_365 = _T_3 ? 8'h0 : _GEN_357; // @[CPU6502.scala 43:17 721:31]
  wire [15:0] _io_memAddr_T = {8'h1,regSP}; // @[Cat.scala 33:92]
  wire [7:0] _regSP_T_1 = regSP - 8'h1; // @[CPU6502.scala 753:26]
  wire [7:0] status = {flagN,flagV,2'h3,flagD,flagI,flagZ,flagC}; // @[Cat.scala 33:92]
  wire [7:0] _regSP_T_5 = regSP + 8'h1; // @[CPU6502.scala 770:28]
  wire [15:0] _GEN_368 = _T_6 ? _io_memAddr_T : regPC; // @[CPU6502.scala 42:14 772:37 773:24]
  wire [7:0] _GEN_374 = _T_3 ? _regSP_T_5 : regSP; // @[CPU6502.scala 769:31 770:19 21:22]
  wire [15:0] _GEN_376 = _T_3 ? regPC : _GEN_368; // @[CPU6502.scala 42:14 769:31]
  wire  _GEN_384 = _T_6 ? io_memDataIn[0] : flagC; // @[CPU6502.scala 786:37 790:19 25:22]
  wire  _GEN_385 = _T_6 ? io_memDataIn[1] : flagZ; // @[CPU6502.scala 786:37 791:19 26:22]
  wire  _GEN_386 = _T_6 ? io_memDataIn[2] : flagI; // @[CPU6502.scala 786:37 792:19 27:22]
  wire  _GEN_387 = _T_6 ? io_memDataIn[3] : flagD; // @[CPU6502.scala 786:37 793:19 28:22]
  wire  _GEN_395 = _T_3 ? flagC : _GEN_384; // @[CPU6502.scala 25:22 783:31]
  wire  _GEN_396 = _T_3 ? flagZ : _GEN_385; // @[CPU6502.scala 26:22 783:31]
  wire  _GEN_397 = _T_3 ? flagI : _GEN_386; // @[CPU6502.scala 27:22 783:31]
  wire  _GEN_398 = _T_3 ? flagD : _GEN_387; // @[CPU6502.scala 28:22 783:31]
  wire  _T_123 = cycle == 3'h3; // @[CPU6502.scala 820:28]
  wire [15:0] _GEN_402 = cycle == 3'h3 ? _io_memAddr_T : regPC; // @[CPU6502.scala 42:14 820:37 822:24]
  wire [7:0] _GEN_403 = cycle == 3'h3 ? regPC[7:0] : 8'h0; // @[CPU6502.scala 43:17 820:37 823:27]
  wire [7:0] _GEN_405 = cycle == 3'h3 ? _regSP_T_1 : regSP; // @[CPU6502.scala 820:37 825:19 21:22]
  wire [15:0] _GEN_406 = cycle == 3'h3 ? operand : regPC; // @[CPU6502.scala 820:37 826:19 22:22]
  wire [1:0] _GEN_407 = cycle == 3'h3 ? 2'h0 : state; // @[CPU6502.scala 820:37 827:19 35:22]
  wire [15:0] _GEN_408 = _T_79 ? _io_memAddr_T : _GEN_402; // @[CPU6502.scala 813:37 815:24]
  wire [7:0] _GEN_409 = _T_79 ? regPC[15:8] : _GEN_403; // @[CPU6502.scala 813:37 816:27]
  wire  _GEN_410 = _T_79 | _T_123; // @[CPU6502.scala 813:37 817:25]
  wire [7:0] _GEN_411 = _T_79 ? _regSP_T_1 : _GEN_405; // @[CPU6502.scala 813:37 818:19]
  wire [2:0] _GEN_412 = _T_79 ? 3'h3 : cycle; // @[CPU6502.scala 813:37 819:19 39:22]
  wire [15:0] _GEN_413 = _T_79 ? regPC : _GEN_406; // @[CPU6502.scala 22:22 813:37]
  wire [1:0] _GEN_414 = _T_79 ? state : _GEN_407; // @[CPU6502.scala 35:22 813:37]
  wire [15:0] _GEN_415 = _T_6 ? regPC : _GEN_408; // @[CPU6502.scala 808:37 809:24]
  wire [15:0] _GEN_417 = _T_6 ? _regPC_T_25 : operand; // @[CPU6502.scala 808:37 811:21 38:24]
  wire [2:0] _GEN_418 = _T_6 ? 3'h2 : _GEN_412; // @[CPU6502.scala 808:37 812:19]
  wire [7:0] _GEN_419 = _T_6 ? 8'h0 : _GEN_409; // @[CPU6502.scala 43:17 808:37]
  wire  _GEN_420 = _T_6 ? 1'h0 : _GEN_410; // @[CPU6502.scala 44:15 808:37]
  wire [7:0] _GEN_421 = _T_6 ? regSP : _GEN_411; // @[CPU6502.scala 21:22 808:37]
  wire [15:0] _GEN_422 = _T_6 ? regPC : _GEN_413; // @[CPU6502.scala 22:22 808:37]
  wire [1:0] _GEN_423 = _T_6 ? state : _GEN_414; // @[CPU6502.scala 35:22 808:37]
  wire [15:0] _GEN_424 = _T_3 ? regPC : _GEN_415; // @[CPU6502.scala 802:31 803:24]
  wire [15:0] _GEN_426 = _T_3 ? {{8'd0}, io_memDataIn} : _GEN_417; // @[CPU6502.scala 802:31 805:21]
  wire [15:0] _GEN_427 = _T_3 ? _regPC_T_1 : _GEN_422; // @[CPU6502.scala 802:31 806:19]
  wire [2:0] _GEN_428 = _T_3 ? 3'h1 : _GEN_418; // @[CPU6502.scala 802:31 807:19]
  wire [7:0] _GEN_429 = _T_3 ? 8'h0 : _GEN_419; // @[CPU6502.scala 43:17 802:31]
  wire  _GEN_430 = _T_3 ? 1'h0 : _GEN_420; // @[CPU6502.scala 44:15 802:31]
  wire [7:0] _GEN_431 = _T_3 ? regSP : _GEN_421; // @[CPU6502.scala 21:22 802:31]
  wire [1:0] _GEN_432 = _T_3 ? state : _GEN_423; // @[CPU6502.scala 35:22 802:31]
  wire [15:0] _regPC_T_113 = _regPC_T_25 + 16'h1; // @[CPU6502.scala 845:55]
  wire [15:0] _GEN_433 = _T_79 ? _io_memAddr_T : regPC; // @[CPU6502.scala 42:14 842:37 843:24]
  wire [15:0] _GEN_435 = _T_79 ? _regPC_T_113 : regPC; // @[CPU6502.scala 842:37 845:19 22:22]
  wire [15:0] _GEN_437 = _T_6 ? _io_memAddr_T : _GEN_433; // @[CPU6502.scala 836:37 837:24]
  wire  _GEN_438 = _T_6 | _T_79; // @[CPU6502.scala 836:37 838:24]
  wire [15:0] _GEN_439 = _T_6 ? {{8'd0}, io_memDataIn} : operand; // @[CPU6502.scala 836:37 839:21 38:24]
  wire [7:0] _GEN_440 = _T_6 ? _regSP_T_5 : regSP; // @[CPU6502.scala 836:37 840:19 21:22]
  wire [15:0] _GEN_442 = _T_6 ? regPC : _GEN_435; // @[CPU6502.scala 22:22 836:37]
  wire [7:0] _GEN_444 = _T_3 ? _regSP_T_5 : _GEN_440; // @[CPU6502.scala 833:31 834:19]
  wire [15:0] _GEN_446 = _T_3 ? regPC : _GEN_437; // @[CPU6502.scala 42:14 833:31]
  wire  _GEN_447 = _T_3 ? 1'h0 : _GEN_438; // @[CPU6502.scala 45:14 833:31]
  wire [15:0] _GEN_448 = _T_3 ? operand : _GEN_439; // @[CPU6502.scala 38:24 833:31]
  wire [15:0] _GEN_449 = _T_3 ? regPC : _GEN_442; // @[CPU6502.scala 22:22 833:31]
  wire  _T_134 = cycle == 3'h5; // @[CPU6502.scala 885:28]
  wire [15:0] _GEN_451 = cycle == 3'h5 ? 16'hffff : regPC; // @[CPU6502.scala 42:14 885:37 887:24]
  wire [15:0] _GEN_453 = cycle == 3'h5 ? _regPC_T_25 : regPC; // @[CPU6502.scala 885:37 889:19 22:22]
  wire [1:0] _GEN_454 = cycle == 3'h5 ? 2'h0 : state; // @[CPU6502.scala 885:37 890:19 35:22]
  wire [15:0] _GEN_455 = cycle == 3'h4 ? 16'hfffe : _GEN_451; // @[CPU6502.scala 879:37 881:24]
  wire  _GEN_456 = cycle == 3'h4 | _T_134; // @[CPU6502.scala 879:37 882:24]
  wire [15:0] _GEN_457 = cycle == 3'h4 ? {{8'd0}, io_memDataIn} : operand; // @[CPU6502.scala 879:37 883:21 38:24]
  wire [2:0] _GEN_458 = cycle == 3'h4 ? 3'h5 : cycle; // @[CPU6502.scala 879:37 884:19 39:22]
  wire [15:0] _GEN_459 = cycle == 3'h4 ? regPC : _GEN_453; // @[CPU6502.scala 22:22 879:37]
  wire [1:0] _GEN_460 = cycle == 3'h4 ? state : _GEN_454; // @[CPU6502.scala 35:22 879:37]
  wire [15:0] _GEN_461 = _T_123 ? _io_memAddr_T : _GEN_455; // @[CPU6502.scala 869:37 872:24]
  wire [7:0] _GEN_462 = _T_123 ? status : 8'h0; // @[CPU6502.scala 43:17 869:37 873:27]
  wire  _GEN_465 = _T_123 | flagI; // @[CPU6502.scala 869:37 876:19 27:22]
  wire [2:0] _GEN_467 = _T_123 ? 3'h4 : _GEN_458; // @[CPU6502.scala 869:37 878:19]
  wire  _GEN_468 = _T_123 ? 1'h0 : _GEN_456; // @[CPU6502.scala 45:14 869:37]
  wire [15:0] _GEN_469 = _T_123 ? operand : _GEN_457; // @[CPU6502.scala 38:24 869:37]
  wire [15:0] _GEN_470 = _T_123 ? regPC : _GEN_459; // @[CPU6502.scala 22:22 869:37]
  wire [1:0] _GEN_471 = _T_123 ? state : _GEN_460; // @[CPU6502.scala 35:22 869:37]
  wire [15:0] _GEN_472 = _T_79 ? _io_memAddr_T : _GEN_461; // @[CPU6502.scala 862:37 864:24]
  wire [7:0] _GEN_473 = _T_79 ? regPC[7:0] : _GEN_462; // @[CPU6502.scala 862:37 865:27]
  wire [2:0] _GEN_476 = _T_79 ? 3'h3 : _GEN_467; // @[CPU6502.scala 862:37 868:19]
  wire  _GEN_477 = _T_79 ? flagI : _GEN_465; // @[CPU6502.scala 27:22 862:37]
  wire  _GEN_479 = _T_79 ? 1'h0 : _GEN_468; // @[CPU6502.scala 45:14 862:37]
  wire [15:0] _GEN_480 = _T_79 ? operand : _GEN_469; // @[CPU6502.scala 38:24 862:37]
  wire [15:0] _GEN_481 = _T_79 ? regPC : _GEN_470; // @[CPU6502.scala 22:22 862:37]
  wire [1:0] _GEN_482 = _T_79 ? state : _GEN_471; // @[CPU6502.scala 35:22 862:37]
  wire [15:0] _GEN_483 = _T_6 ? _io_memAddr_T : _GEN_472; // @[CPU6502.scala 855:37 857:24]
  wire [7:0] _GEN_484 = _T_6 ? regPC[15:8] : _GEN_473; // @[CPU6502.scala 855:37 858:27]
  wire  _GEN_485 = _T_6 | _GEN_410; // @[CPU6502.scala 855:37 859:25]
  wire [7:0] _GEN_486 = _T_6 ? _regSP_T_1 : _GEN_411; // @[CPU6502.scala 855:37 860:19]
  wire [2:0] _GEN_487 = _T_6 ? 3'h2 : _GEN_476; // @[CPU6502.scala 855:37 861:19]
  wire  _GEN_488 = _T_6 ? flagI : _GEN_477; // @[CPU6502.scala 27:22 855:37]
  wire  _GEN_490 = _T_6 ? 1'h0 : _GEN_479; // @[CPU6502.scala 45:14 855:37]
  wire [15:0] _GEN_491 = _T_6 ? operand : _GEN_480; // @[CPU6502.scala 38:24 855:37]
  wire [15:0] _GEN_492 = _T_6 ? regPC : _GEN_481; // @[CPU6502.scala 22:22 855:37]
  wire [1:0] _GEN_493 = _T_6 ? state : _GEN_482; // @[CPU6502.scala 35:22 855:37]
  wire [15:0] _GEN_494 = _T_3 ? _regPC_T_1 : _GEN_492; // @[CPU6502.scala 852:31 853:19]
  wire [2:0] _GEN_495 = _T_3 ? 3'h1 : _GEN_487; // @[CPU6502.scala 852:31 854:19]
  wire [15:0] _GEN_496 = _T_3 ? regPC : _GEN_483; // @[CPU6502.scala 42:14 852:31]
  wire [7:0] _GEN_497 = _T_3 ? 8'h0 : _GEN_484; // @[CPU6502.scala 43:17 852:31]
  wire  _GEN_498 = _T_3 ? 1'h0 : _GEN_485; // @[CPU6502.scala 44:15 852:31]
  wire [7:0] _GEN_499 = _T_3 ? regSP : _GEN_486; // @[CPU6502.scala 21:22 852:31]
  wire  _GEN_500 = _T_3 ? flagI : _GEN_488; // @[CPU6502.scala 27:22 852:31]
  wire  _GEN_502 = _T_3 ? 1'h0 : _GEN_490; // @[CPU6502.scala 45:14 852:31]
  wire [15:0] _GEN_503 = _T_3 ? operand : _GEN_491; // @[CPU6502.scala 38:24 852:31]
  wire [1:0] _GEN_504 = _T_3 ? state : _GEN_493; // @[CPU6502.scala 35:22 852:31]
  wire [15:0] _GEN_507 = _T_123 ? _regPC_T_25 : regPC; // @[CPU6502.scala 919:37 923:19 22:22]
  wire [15:0] _GEN_511 = _T_79 ? {{8'd0}, io_memDataIn} : operand; // @[CPU6502.scala 912:37 916:21 38:24]
  wire [7:0] _GEN_512 = _T_79 ? _regSP_T_5 : regSP; // @[CPU6502.scala 912:37 917:19 21:22]
  wire [15:0] _GEN_514 = _T_79 ? regPC : _GEN_507; // @[CPU6502.scala 22:22 912:37]
  wire [15:0] _GEN_516 = _T_6 ? _io_memAddr_T : _GEN_408; // @[CPU6502.scala 899:37 901:24]
  wire [7:0] _GEN_524 = _T_6 ? _regSP_T_5 : _GEN_512; // @[CPU6502.scala 899:37 910:19]
  wire [15:0] _GEN_526 = _T_6 ? operand : _GEN_511; // @[CPU6502.scala 38:24 899:37]
  wire [15:0] _GEN_527 = _T_6 ? regPC : _GEN_514; // @[CPU6502.scala 22:22 899:37]
  wire [7:0] _GEN_529 = _T_3 ? _regSP_T_5 : _GEN_524; // @[CPU6502.scala 896:31 897:19]
  wire [15:0] _GEN_531 = _T_3 ? regPC : _GEN_516; // @[CPU6502.scala 42:14 896:31]
  wire [15:0] _GEN_539 = _T_3 ? operand : _GEN_526; // @[CPU6502.scala 38:24 896:31]
  wire [15:0] _GEN_540 = _T_3 ? regPC : _GEN_527; // @[CPU6502.scala 22:22 896:31]
  wire [7:0] _GEN_544 = _T_79 ? io_memDataIn : regA; // @[CPU6502.scala 942:37 945:18 18:21]
  wire  _GEN_545 = _T_79 ? io_memDataIn[7] : flagN; // @[CPU6502.scala 50:11 31:22 942:37]
  wire  _GEN_546 = _T_79 ? io_memDataIn == 8'h0 : flagZ; // @[CPU6502.scala 51:11 26:22 942:37]
  wire [15:0] _GEN_548 = _T_6 ? regPC : _GEN_188; // @[CPU6502.scala 936:37 937:24]
  wire [15:0] _GEN_551 = _T_6 ? _regPC_T_1 : regPC; // @[CPU6502.scala 936:37 940:19 22:22]
  wire [7:0] _GEN_553 = _T_6 ? regA : _GEN_544; // @[CPU6502.scala 18:21 936:37]
  wire  _GEN_554 = _T_6 ? flagN : _GEN_545; // @[CPU6502.scala 31:22 936:37]
  wire  _GEN_555 = _T_6 ? flagZ : _GEN_546; // @[CPU6502.scala 26:22 936:37]
  wire [15:0] _GEN_557 = _T_3 ? regPC : _GEN_548; // @[CPU6502.scala 930:31 931:24]
  wire  _GEN_558 = _T_3 | _GEN_438; // @[CPU6502.scala 930:31 932:24]
  wire [15:0] _GEN_560 = _T_3 ? _regPC_T_1 : _GEN_551; // @[CPU6502.scala 930:31 934:19]
  wire [7:0] _GEN_562 = _T_3 ? regA : _GEN_553; // @[CPU6502.scala 18:21 930:31]
  wire  _GEN_563 = _T_3 ? flagN : _GEN_554; // @[CPU6502.scala 31:22 930:31]
  wire  _GEN_564 = _T_3 ? flagZ : _GEN_555; // @[CPU6502.scala 26:22 930:31]
  wire [7:0] _GEN_567 = _T_79 ? regA : 8'h0; // @[CPU6502.scala 43:17 965:37 967:27]
  wire [7:0] _GEN_575 = _T_6 ? 8'h0 : _GEN_567; // @[CPU6502.scala 43:17 959:37]
  wire [7:0] _GEN_583 = _T_3 ? 8'h0 : _GEN_575; // @[CPU6502.scala 43:17 953:31]
  wire [7:0] _operand_T_7 = io_memDataIn + regX; // @[CPU6502.scala 978:52]
  wire [15:0] _operand_T_9 = {8'h0,_operand_T_7}; // @[Cat.scala 33:92]
  wire [15:0] _GEN_594 = _T_3 ? _operand_T_9 : operand; // @[CPU6502.scala 975:31 978:21 38:24]
  wire [15:0] _GEN_1902 = {{8'd0}, regX}; // @[CPU6502.scala 1017:57]
  wire [15:0] _operand_T_17 = _regPC_T_25 + _GEN_1902; // @[CPU6502.scala 1017:57]
  wire [15:0] _GEN_621 = _T_6 ? _operand_T_17 : operand; // @[CPU6502.scala 1014:37 1017:21 38:24]
  wire [15:0] _GEN_630 = _T_3 ? {{8'd0}, io_memDataIn} : _GEN_621; // @[CPU6502.scala 1008:31 1011:21]
  wire [15:0] _GEN_1903 = {{8'd0}, regY}; // @[CPU6502.scala 1040:57]
  wire [15:0] _operand_T_21 = _regPC_T_25 + _GEN_1903; // @[CPU6502.scala 1040:57]
  wire [15:0] _GEN_645 = _T_6 ? _operand_T_21 : operand; // @[CPU6502.scala 1037:37 1040:21 38:24]
  wire [15:0] _GEN_654 = _T_3 ? {{8'd0}, io_memDataIn} : _GEN_645; // @[CPU6502.scala 1031:31 1034:21]
  wire [7:0] result_21 = regA + 8'h1; // @[CPU6502.scala 1054:29]
  wire [7:0] result_22 = regA - 8'h1; // @[CPU6502.scala 1062:29]
  wire [7:0] _GEN_661 = 8'h3a == opcode ? result_22 : regA; // @[CPU6502.scala 1063:16 18:21 66:22]
  wire  _GEN_662 = 8'h3a == opcode ? result_22[7] : flagN; // @[CPU6502.scala 50:11 31:22 66:22]
  wire  _GEN_663 = 8'h3a == opcode ? result_22 == 8'h0 : flagZ; // @[CPU6502.scala 51:11 26:22 66:22]
  wire [1:0] _GEN_664 = 8'h3a == opcode ? 2'h0 : state; // @[CPU6502.scala 1065:17 35:22 66:22]
  wire [7:0] _GEN_665 = 8'h1a == opcode ? result_21 : _GEN_661; // @[CPU6502.scala 1055:16 66:22]
  wire  _GEN_666 = 8'h1a == opcode ? result_21[7] : _GEN_662; // @[CPU6502.scala 50:11 66:22]
  wire  _GEN_667 = 8'h1a == opcode ? result_21 == 8'h0 : _GEN_663; // @[CPU6502.scala 51:11 66:22]
  wire [1:0] _GEN_668 = 8'h1a == opcode ? 2'h0 : _GEN_664; // @[CPU6502.scala 1057:17 66:22]
  wire [15:0] _GEN_669 = 8'hb9 == opcode ? _GEN_557 : regPC; // @[CPU6502.scala 42:14 66:22]
  wire  _GEN_670 = 8'hb9 == opcode & _GEN_558; // @[CPU6502.scala 45:14 66:22]
  wire [15:0] _GEN_671 = 8'hb9 == opcode ? _GEN_654 : operand; // @[CPU6502.scala 66:22 38:24]
  wire [15:0] _GEN_672 = 8'hb9 == opcode ? _GEN_560 : regPC; // @[CPU6502.scala 22:22 66:22]
  wire [2:0] _GEN_673 = 8'hb9 == opcode ? _GEN_208 : cycle; // @[CPU6502.scala 39:22 66:22]
  wire [7:0] _GEN_674 = 8'hb9 == opcode ? _GEN_562 : _GEN_665; // @[CPU6502.scala 66:22]
  wire  _GEN_675 = 8'hb9 == opcode ? _GEN_563 : _GEN_666; // @[CPU6502.scala 66:22]
  wire  _GEN_676 = 8'hb9 == opcode ? _GEN_564 : _GEN_667; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_677 = 8'hb9 == opcode ? _GEN_214 : _GEN_668; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_678 = 8'hbd == opcode ? _GEN_557 : _GEN_669; // @[CPU6502.scala 66:22]
  wire  _GEN_679 = 8'hbd == opcode ? _GEN_558 : _GEN_670; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_680 = 8'hbd == opcode ? _GEN_630 : _GEN_671; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_681 = 8'hbd == opcode ? _GEN_560 : _GEN_672; // @[CPU6502.scala 66:22]
  wire [2:0] _GEN_682 = 8'hbd == opcode ? _GEN_208 : _GEN_673; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_683 = 8'hbd == opcode ? _GEN_562 : _GEN_674; // @[CPU6502.scala 66:22]
  wire  _GEN_684 = 8'hbd == opcode ? _GEN_563 : _GEN_675; // @[CPU6502.scala 66:22]
  wire  _GEN_685 = 8'hbd == opcode ? _GEN_564 : _GEN_676; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_686 = 8'hbd == opcode ? _GEN_214 : _GEN_677; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_687 = 8'h95 == opcode ? _GEN_13 : _GEN_678; // @[CPU6502.scala 66:22]
  wire  _GEN_688 = 8'h95 == opcode ? _T_3 : _GEN_679; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_689 = 8'h95 == opcode ? _GEN_594 : _GEN_680; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_690 = 8'h95 == opcode ? _GEN_5 : _GEN_681; // @[CPU6502.scala 66:22]
  wire [2:0] _GEN_691 = 8'h95 == opcode ? _GEN_17 : _GEN_682; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_692 = 8'h95 == opcode ? _GEN_45 : 8'h0; // @[CPU6502.scala 43:17 66:22]
  wire [1:0] _GEN_694 = 8'h95 == opcode ? _GEN_21 : _GEN_686; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_695 = 8'h95 == opcode ? regA : _GEN_683; // @[CPU6502.scala 18:21 66:22]
  wire  _GEN_696 = 8'h95 == opcode ? flagN : _GEN_684; // @[CPU6502.scala 31:22 66:22]
  wire  _GEN_697 = 8'h95 == opcode ? flagZ : _GEN_685; // @[CPU6502.scala 26:22 66:22]
  wire [15:0] _GEN_698 = 8'hb5 == opcode ? _GEN_13 : _GEN_687; // @[CPU6502.scala 66:22]
  wire  _GEN_699 = 8'hb5 == opcode ? _GEN_14 : _GEN_688; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_700 = 8'hb5 == opcode ? _GEN_594 : _GEN_689; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_701 = 8'hb5 == opcode ? _GEN_5 : _GEN_690; // @[CPU6502.scala 66:22]
  wire [2:0] _GEN_702 = 8'hb5 == opcode ? _GEN_17 : _GEN_691; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_703 = 8'hb5 == opcode ? _GEN_18 : _GEN_695; // @[CPU6502.scala 66:22]
  wire  _GEN_704 = 8'hb5 == opcode ? _GEN_19 : _GEN_696; // @[CPU6502.scala 66:22]
  wire  _GEN_705 = 8'hb5 == opcode ? _GEN_20 : _GEN_697; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_706 = 8'hb5 == opcode ? _GEN_21 : _GEN_694; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_707 = 8'hb5 == opcode ? 8'h0 : _GEN_692; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_708 = 8'hb5 == opcode ? 1'h0 : 8'h95 == opcode & _GEN_46; // @[CPU6502.scala 44:15 66:22]
  wire [15:0] _GEN_709 = 8'h8d == opcode ? _GEN_557 : _GEN_698; // @[CPU6502.scala 66:22]
  wire  _GEN_710 = 8'h8d == opcode ? _GEN_14 : _GEN_699; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_711 = 8'h8d == opcode ? _GEN_426 : _GEN_700; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_712 = 8'h8d == opcode ? _GEN_560 : _GEN_701; // @[CPU6502.scala 66:22]
  wire [2:0] _GEN_713 = 8'h8d == opcode ? _GEN_208 : _GEN_702; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_714 = 8'h8d == opcode ? _GEN_583 : _GEN_707; // @[CPU6502.scala 66:22]
  wire  _GEN_715 = 8'h8d == opcode ? _GEN_211 : _GEN_708; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_716 = 8'h8d == opcode ? _GEN_214 : _GEN_706; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_717 = 8'h8d == opcode ? regA : _GEN_703; // @[CPU6502.scala 18:21 66:22]
  wire  _GEN_718 = 8'h8d == opcode ? flagN : _GEN_704; // @[CPU6502.scala 31:22 66:22]
  wire  _GEN_719 = 8'h8d == opcode ? flagZ : _GEN_705; // @[CPU6502.scala 26:22 66:22]
  wire [15:0] _GEN_720 = 8'had == opcode ? _GEN_557 : _GEN_709; // @[CPU6502.scala 66:22]
  wire  _GEN_721 = 8'had == opcode ? _GEN_558 : _GEN_710; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_722 = 8'had == opcode ? _GEN_426 : _GEN_711; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_723 = 8'had == opcode ? _GEN_560 : _GEN_712; // @[CPU6502.scala 66:22]
  wire [2:0] _GEN_724 = 8'had == opcode ? _GEN_208 : _GEN_713; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_725 = 8'had == opcode ? _GEN_562 : _GEN_717; // @[CPU6502.scala 66:22]
  wire  _GEN_726 = 8'had == opcode ? _GEN_563 : _GEN_718; // @[CPU6502.scala 66:22]
  wire  _GEN_727 = 8'had == opcode ? _GEN_564 : _GEN_719; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_728 = 8'had == opcode ? _GEN_214 : _GEN_716; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_729 = 8'had == opcode ? 8'h0 : _GEN_714; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_730 = 8'had == opcode ? 1'h0 : _GEN_715; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_731 = 8'h40 == opcode ? _GEN_529 : regSP; // @[CPU6502.scala 21:22 66:22]
  wire [2:0] _GEN_732 = 8'h40 == opcode ? _GEN_428 : _GEN_724; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_733 = 8'h40 == opcode ? _GEN_531 : _GEN_720; // @[CPU6502.scala 66:22]
  wire  _GEN_734 = 8'h40 == opcode ? _GEN_498 : _GEN_721; // @[CPU6502.scala 66:22]
  wire  _GEN_735 = 8'h40 == opcode ? _GEN_395 : flagC; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_736 = 8'h40 == opcode ? _GEN_396 : _GEN_727; // @[CPU6502.scala 66:22]
  wire  _GEN_737 = 8'h40 == opcode ? _GEN_397 : flagI; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_738 = 8'h40 == opcode ? _GEN_398 : flagD; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_739 = 8'h40 == opcode ? _GEN_186 : flagV; // @[CPU6502.scala 30:22 66:22]
  wire  _GEN_740 = 8'h40 == opcode ? _GEN_19 : _GEN_726; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_741 = 8'h40 == opcode ? _GEN_539 : _GEN_722; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_742 = 8'h40 == opcode ? _GEN_540 : _GEN_723; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_743 = 8'h40 == opcode ? _GEN_432 : _GEN_728; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_744 = 8'h40 == opcode ? regA : _GEN_725; // @[CPU6502.scala 18:21 66:22]
  wire [7:0] _GEN_745 = 8'h40 == opcode ? 8'h0 : _GEN_729; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_746 = 8'h40 == opcode ? 1'h0 : _GEN_730; // @[CPU6502.scala 44:15 66:22]
  wire [15:0] _GEN_747 = 8'h0 == opcode ? _GEN_494 : _GEN_742; // @[CPU6502.scala 66:22]
  wire [2:0] _GEN_748 = 8'h0 == opcode ? _GEN_495 : _GEN_732; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_749 = 8'h0 == opcode ? _GEN_496 : _GEN_733; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_750 = 8'h0 == opcode ? _GEN_497 : _GEN_745; // @[CPU6502.scala 66:22]
  wire  _GEN_751 = 8'h0 == opcode ? _GEN_498 : _GEN_746; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_752 = 8'h0 == opcode ? _GEN_499 : _GEN_731; // @[CPU6502.scala 66:22]
  wire  _GEN_753 = 8'h0 == opcode ? _GEN_500 : _GEN_737; // @[CPU6502.scala 66:22]
  wire  _GEN_755 = 8'h0 == opcode ? _GEN_502 : _GEN_734; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_756 = 8'h0 == opcode ? _GEN_503 : _GEN_741; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_757 = 8'h0 == opcode ? _GEN_504 : _GEN_743; // @[CPU6502.scala 66:22]
  wire  _GEN_758 = 8'h0 == opcode ? flagC : _GEN_735; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_759 = 8'h0 == opcode ? flagZ : _GEN_736; // @[CPU6502.scala 26:22 66:22]
  wire  _GEN_760 = 8'h0 == opcode ? flagD : _GEN_738; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_761 = 8'h0 == opcode ? flagV : _GEN_739; // @[CPU6502.scala 30:22 66:22]
  wire  _GEN_762 = 8'h0 == opcode ? flagN : _GEN_740; // @[CPU6502.scala 31:22 66:22]
  wire [7:0] _GEN_763 = 8'h0 == opcode ? regA : _GEN_744; // @[CPU6502.scala 18:21 66:22]
  wire [7:0] _GEN_764 = 8'h60 == opcode ? _GEN_444 : _GEN_752; // @[CPU6502.scala 66:22]
  wire [2:0] _GEN_765 = 8'h60 == opcode ? _GEN_208 : _GEN_748; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_766 = 8'h60 == opcode ? _GEN_446 : _GEN_749; // @[CPU6502.scala 66:22]
  wire  _GEN_767 = 8'h60 == opcode ? _GEN_447 : _GEN_755; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_768 = 8'h60 == opcode ? _GEN_448 : _GEN_756; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_769 = 8'h60 == opcode ? _GEN_449 : _GEN_747; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_770 = 8'h60 == opcode ? _GEN_214 : _GEN_757; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_771 = 8'h60 == opcode ? 8'h0 : _GEN_750; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_772 = 8'h60 == opcode ? 1'h0 : _GEN_751; // @[CPU6502.scala 44:15 66:22]
  wire  _GEN_773 = 8'h60 == opcode ? flagI : _GEN_753; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_775 = 8'h60 == opcode ? flagC : _GEN_758; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_776 = 8'h60 == opcode ? flagZ : _GEN_759; // @[CPU6502.scala 26:22 66:22]
  wire  _GEN_777 = 8'h60 == opcode ? flagD : _GEN_760; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_778 = 8'h60 == opcode ? flagV : _GEN_761; // @[CPU6502.scala 30:22 66:22]
  wire  _GEN_779 = 8'h60 == opcode ? flagN : _GEN_762; // @[CPU6502.scala 31:22 66:22]
  wire [7:0] _GEN_780 = 8'h60 == opcode ? regA : _GEN_763; // @[CPU6502.scala 18:21 66:22]
  wire [15:0] _GEN_781 = 8'h20 == opcode ? _GEN_424 : _GEN_766; // @[CPU6502.scala 66:22]
  wire  _GEN_782 = 8'h20 == opcode ? _GEN_14 : _GEN_767; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_783 = 8'h20 == opcode ? _GEN_426 : _GEN_768; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_784 = 8'h20 == opcode ? _GEN_427 : _GEN_769; // @[CPU6502.scala 66:22]
  wire [2:0] _GEN_785 = 8'h20 == opcode ? _GEN_428 : _GEN_765; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_786 = 8'h20 == opcode ? _GEN_429 : _GEN_771; // @[CPU6502.scala 66:22]
  wire  _GEN_787 = 8'h20 == opcode ? _GEN_430 : _GEN_772; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_788 = 8'h20 == opcode ? _GEN_431 : _GEN_764; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_789 = 8'h20 == opcode ? _GEN_432 : _GEN_770; // @[CPU6502.scala 66:22]
  wire  _GEN_790 = 8'h20 == opcode ? flagI : _GEN_773; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_792 = 8'h20 == opcode ? flagC : _GEN_775; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_793 = 8'h20 == opcode ? flagZ : _GEN_776; // @[CPU6502.scala 26:22 66:22]
  wire  _GEN_794 = 8'h20 == opcode ? flagD : _GEN_777; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_795 = 8'h20 == opcode ? flagV : _GEN_778; // @[CPU6502.scala 30:22 66:22]
  wire  _GEN_796 = 8'h20 == opcode ? flagN : _GEN_779; // @[CPU6502.scala 31:22 66:22]
  wire [7:0] _GEN_797 = 8'h20 == opcode ? regA : _GEN_780; // @[CPU6502.scala 18:21 66:22]
  wire [7:0] _GEN_798 = 8'h28 == opcode ? _GEN_374 : _GEN_788; // @[CPU6502.scala 66:22]
  wire [2:0] _GEN_799 = 8'h28 == opcode ? _GEN_17 : _GEN_785; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_800 = 8'h28 == opcode ? _GEN_376 : _GEN_781; // @[CPU6502.scala 66:22]
  wire  _GEN_801 = 8'h28 == opcode ? _GEN_46 : _GEN_782; // @[CPU6502.scala 66:22]
  wire  _GEN_802 = 8'h28 == opcode ? _GEN_395 : _GEN_792; // @[CPU6502.scala 66:22]
  wire  _GEN_803 = 8'h28 == opcode ? _GEN_396 : _GEN_793; // @[CPU6502.scala 66:22]
  wire  _GEN_804 = 8'h28 == opcode ? _GEN_397 : _GEN_790; // @[CPU6502.scala 66:22]
  wire  _GEN_805 = 8'h28 == opcode ? _GEN_398 : _GEN_794; // @[CPU6502.scala 66:22]
  wire  _GEN_806 = 8'h28 == opcode ? _GEN_186 : _GEN_795; // @[CPU6502.scala 66:22]
  wire  _GEN_807 = 8'h28 == opcode ? _GEN_19 : _GEN_796; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_808 = 8'h28 == opcode ? _GEN_21 : _GEN_789; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_809 = 8'h28 == opcode ? operand : _GEN_783; // @[CPU6502.scala 66:22 38:24]
  wire [15:0] _GEN_810 = 8'h28 == opcode ? regPC : _GEN_784; // @[CPU6502.scala 22:22 66:22]
  wire [7:0] _GEN_811 = 8'h28 == opcode ? 8'h0 : _GEN_786; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_812 = 8'h28 == opcode ? 1'h0 : _GEN_787; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_814 = 8'h28 == opcode ? regA : _GEN_797; // @[CPU6502.scala 18:21 66:22]
  wire [7:0] _GEN_815 = 8'h68 == opcode ? _GEN_374 : _GEN_798; // @[CPU6502.scala 66:22]
  wire [2:0] _GEN_816 = 8'h68 == opcode ? _GEN_17 : _GEN_799; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_817 = 8'h68 == opcode ? _GEN_376 : _GEN_800; // @[CPU6502.scala 66:22]
  wire  _GEN_818 = 8'h68 == opcode ? _GEN_46 : _GEN_801; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_819 = 8'h68 == opcode ? _GEN_18 : _GEN_814; // @[CPU6502.scala 66:22]
  wire  _GEN_820 = 8'h68 == opcode ? _GEN_19 : _GEN_807; // @[CPU6502.scala 66:22]
  wire  _GEN_821 = 8'h68 == opcode ? _GEN_20 : _GEN_803; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_822 = 8'h68 == opcode ? _GEN_21 : _GEN_808; // @[CPU6502.scala 66:22]
  wire  _GEN_823 = 8'h68 == opcode ? flagC : _GEN_802; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_824 = 8'h68 == opcode ? flagI : _GEN_804; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_825 = 8'h68 == opcode ? flagD : _GEN_805; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_826 = 8'h68 == opcode ? flagV : _GEN_806; // @[CPU6502.scala 30:22 66:22]
  wire [15:0] _GEN_827 = 8'h68 == opcode ? operand : _GEN_809; // @[CPU6502.scala 66:22 38:24]
  wire [15:0] _GEN_828 = 8'h68 == opcode ? regPC : _GEN_810; // @[CPU6502.scala 22:22 66:22]
  wire [7:0] _GEN_829 = 8'h68 == opcode ? 8'h0 : _GEN_811; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_830 = 8'h68 == opcode ? 1'h0 : _GEN_812; // @[CPU6502.scala 44:15 66:22]
  wire [15:0] _GEN_832 = 8'h8 == opcode ? _io_memAddr_T : _GEN_817; // @[CPU6502.scala 66:22 760:22]
  wire [7:0] _GEN_833 = 8'h8 == opcode ? status : _GEN_829; // @[CPU6502.scala 66:22 761:25]
  wire  _GEN_834 = 8'h8 == opcode | _GEN_830; // @[CPU6502.scala 66:22 762:23]
  wire [7:0] _GEN_835 = 8'h8 == opcode ? _regSP_T_1 : _GEN_815; // @[CPU6502.scala 66:22 763:17]
  wire [1:0] _GEN_836 = 8'h8 == opcode ? 2'h0 : _GEN_822; // @[CPU6502.scala 66:22 764:17]
  wire [2:0] _GEN_837 = 8'h8 == opcode ? cycle : _GEN_816; // @[CPU6502.scala 39:22 66:22]
  wire  _GEN_838 = 8'h8 == opcode ? 1'h0 : _GEN_818; // @[CPU6502.scala 45:14 66:22]
  wire [7:0] _GEN_839 = 8'h8 == opcode ? regA : _GEN_819; // @[CPU6502.scala 18:21 66:22]
  wire  _GEN_840 = 8'h8 == opcode ? flagN : _GEN_820; // @[CPU6502.scala 31:22 66:22]
  wire  _GEN_841 = 8'h8 == opcode ? flagZ : _GEN_821; // @[CPU6502.scala 26:22 66:22]
  wire  _GEN_842 = 8'h8 == opcode ? flagC : _GEN_823; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_843 = 8'h8 == opcode ? flagI : _GEN_824; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_844 = 8'h8 == opcode ? flagD : _GEN_825; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_845 = 8'h8 == opcode ? flagV : _GEN_826; // @[CPU6502.scala 30:22 66:22]
  wire [15:0] _GEN_846 = 8'h8 == opcode ? operand : _GEN_827; // @[CPU6502.scala 66:22 38:24]
  wire [15:0] _GEN_847 = 8'h8 == opcode ? regPC : _GEN_828; // @[CPU6502.scala 22:22 66:22]
  wire [15:0] _GEN_849 = 8'h48 == opcode ? _io_memAddr_T : _GEN_832; // @[CPU6502.scala 66:22 750:22]
  wire [7:0] _GEN_850 = 8'h48 == opcode ? regA : _GEN_833; // @[CPU6502.scala 66:22 751:25]
  wire  _GEN_851 = 8'h48 == opcode | _GEN_834; // @[CPU6502.scala 66:22 752:23]
  wire [7:0] _GEN_852 = 8'h48 == opcode ? _regSP_T_1 : _GEN_835; // @[CPU6502.scala 66:22 753:17]
  wire [1:0] _GEN_853 = 8'h48 == opcode ? 2'h0 : _GEN_836; // @[CPU6502.scala 66:22 754:17]
  wire [2:0] _GEN_854 = 8'h48 == opcode ? cycle : _GEN_837; // @[CPU6502.scala 39:22 66:22]
  wire  _GEN_855 = 8'h48 == opcode ? 1'h0 : _GEN_838; // @[CPU6502.scala 45:14 66:22]
  wire [7:0] _GEN_856 = 8'h48 == opcode ? regA : _GEN_839; // @[CPU6502.scala 18:21 66:22]
  wire  _GEN_857 = 8'h48 == opcode ? flagN : _GEN_840; // @[CPU6502.scala 31:22 66:22]
  wire  _GEN_858 = 8'h48 == opcode ? flagZ : _GEN_841; // @[CPU6502.scala 26:22 66:22]
  wire  _GEN_859 = 8'h48 == opcode ? flagC : _GEN_842; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_860 = 8'h48 == opcode ? flagI : _GEN_843; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_861 = 8'h48 == opcode ? flagD : _GEN_844; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_862 = 8'h48 == opcode ? flagV : _GEN_845; // @[CPU6502.scala 30:22 66:22]
  wire [15:0] _GEN_863 = 8'h48 == opcode ? operand : _GEN_846; // @[CPU6502.scala 66:22 38:24]
  wire [15:0] _GEN_864 = 8'h48 == opcode ? regPC : _GEN_847; // @[CPU6502.scala 22:22 66:22]
  wire [7:0] _GEN_866 = 8'h9a == opcode ? regX : _GEN_852; // @[CPU6502.scala 66:22 744:17]
  wire [1:0] _GEN_867 = 8'h9a == opcode ? 2'h0 : _GEN_853; // @[CPU6502.scala 66:22 745:17]
  wire [15:0] _GEN_868 = 8'h9a == opcode ? regPC : _GEN_849; // @[CPU6502.scala 42:14 66:22]
  wire [7:0] _GEN_869 = 8'h9a == opcode ? 8'h0 : _GEN_850; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_870 = 8'h9a == opcode ? 1'h0 : _GEN_851; // @[CPU6502.scala 44:15 66:22]
  wire [2:0] _GEN_871 = 8'h9a == opcode ? cycle : _GEN_854; // @[CPU6502.scala 39:22 66:22]
  wire  _GEN_872 = 8'h9a == opcode ? 1'h0 : _GEN_855; // @[CPU6502.scala 45:14 66:22]
  wire [7:0] _GEN_873 = 8'h9a == opcode ? regA : _GEN_856; // @[CPU6502.scala 18:21 66:22]
  wire  _GEN_874 = 8'h9a == opcode ? flagN : _GEN_857; // @[CPU6502.scala 31:22 66:22]
  wire  _GEN_875 = 8'h9a == opcode ? flagZ : _GEN_858; // @[CPU6502.scala 26:22 66:22]
  wire  _GEN_876 = 8'h9a == opcode ? flagC : _GEN_859; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_877 = 8'h9a == opcode ? flagI : _GEN_860; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_878 = 8'h9a == opcode ? flagD : _GEN_861; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_879 = 8'h9a == opcode ? flagV : _GEN_862; // @[CPU6502.scala 30:22 66:22]
  wire [15:0] _GEN_880 = 8'h9a == opcode ? operand : _GEN_863; // @[CPU6502.scala 66:22 38:24]
  wire [15:0] _GEN_881 = 8'h9a == opcode ? regPC : _GEN_864; // @[CPU6502.scala 22:22 66:22]
  wire [7:0] _GEN_883 = 8'hba == opcode ? regSP : regX; // @[CPU6502.scala 66:22 737:16 19:21]
  wire  _GEN_884 = 8'hba == opcode ? regSP[7] : _GEN_874; // @[CPU6502.scala 50:11 66:22]
  wire  _GEN_885 = 8'hba == opcode ? regSP == 8'h0 : _GEN_875; // @[CPU6502.scala 51:11 66:22]
  wire [1:0] _GEN_886 = 8'hba == opcode ? 2'h0 : _GEN_867; // @[CPU6502.scala 66:22 739:17]
  wire [7:0] _GEN_887 = 8'hba == opcode ? regSP : _GEN_866; // @[CPU6502.scala 21:22 66:22]
  wire [15:0] _GEN_888 = 8'hba == opcode ? regPC : _GEN_868; // @[CPU6502.scala 42:14 66:22]
  wire [7:0] _GEN_889 = 8'hba == opcode ? 8'h0 : _GEN_869; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_890 = 8'hba == opcode ? 1'h0 : _GEN_870; // @[CPU6502.scala 44:15 66:22]
  wire [2:0] _GEN_891 = 8'hba == opcode ? cycle : _GEN_871; // @[CPU6502.scala 39:22 66:22]
  wire  _GEN_892 = 8'hba == opcode ? 1'h0 : _GEN_872; // @[CPU6502.scala 45:14 66:22]
  wire [7:0] _GEN_893 = 8'hba == opcode ? regA : _GEN_873; // @[CPU6502.scala 18:21 66:22]
  wire  _GEN_894 = 8'hba == opcode ? flagC : _GEN_876; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_895 = 8'hba == opcode ? flagI : _GEN_877; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_896 = 8'hba == opcode ? flagD : _GEN_878; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_897 = 8'hba == opcode ? flagV : _GEN_879; // @[CPU6502.scala 30:22 66:22]
  wire [15:0] _GEN_898 = 8'hba == opcode ? operand : _GEN_880; // @[CPU6502.scala 66:22 38:24]
  wire [15:0] _GEN_899 = 8'hba == opcode ? regPC : _GEN_881; // @[CPU6502.scala 22:22 66:22]
  wire [15:0] _GEN_901 = 8'h84 == opcode ? _GEN_13 : _GEN_888; // @[CPU6502.scala 66:22]
  wire  _GEN_902 = 8'h84 == opcode ? _T_3 : _GEN_892; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_903 = 8'h84 == opcode ? _GEN_15 : _GEN_898; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_904 = 8'h84 == opcode ? _GEN_5 : _GEN_899; // @[CPU6502.scala 66:22]
  wire [2:0] _GEN_905 = 8'h84 == opcode ? _GEN_17 : _GEN_891; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_906 = 8'h84 == opcode ? _GEN_365 : _GEN_889; // @[CPU6502.scala 66:22]
  wire  _GEN_907 = 8'h84 == opcode ? _GEN_46 : _GEN_890; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_908 = 8'h84 == opcode ? _GEN_21 : _GEN_886; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_909 = 8'h84 == opcode ? regX : _GEN_883; // @[CPU6502.scala 19:21 66:22]
  wire  _GEN_910 = 8'h84 == opcode ? flagN : _GEN_884; // @[CPU6502.scala 31:22 66:22]
  wire  _GEN_911 = 8'h84 == opcode ? flagZ : _GEN_885; // @[CPU6502.scala 26:22 66:22]
  wire [7:0] _GEN_912 = 8'h84 == opcode ? regSP : _GEN_887; // @[CPU6502.scala 21:22 66:22]
  wire [7:0] _GEN_913 = 8'h84 == opcode ? regA : _GEN_893; // @[CPU6502.scala 18:21 66:22]
  wire  _GEN_914 = 8'h84 == opcode ? flagC : _GEN_894; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_915 = 8'h84 == opcode ? flagI : _GEN_895; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_916 = 8'h84 == opcode ? flagD : _GEN_896; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_917 = 8'h84 == opcode ? flagV : _GEN_897; // @[CPU6502.scala 30:22 66:22]
  wire [15:0] _GEN_919 = 8'h86 == opcode ? _GEN_13 : _GEN_901; // @[CPU6502.scala 66:22]
  wire  _GEN_920 = 8'h86 == opcode ? _T_3 : _GEN_902; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_921 = 8'h86 == opcode ? _GEN_15 : _GEN_903; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_922 = 8'h86 == opcode ? _GEN_5 : _GEN_904; // @[CPU6502.scala 66:22]
  wire [2:0] _GEN_923 = 8'h86 == opcode ? _GEN_17 : _GEN_905; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_924 = 8'h86 == opcode ? _GEN_353 : _GEN_906; // @[CPU6502.scala 66:22]
  wire  _GEN_925 = 8'h86 == opcode ? _GEN_46 : _GEN_907; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_926 = 8'h86 == opcode ? _GEN_21 : _GEN_908; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_927 = 8'h86 == opcode ? regX : _GEN_909; // @[CPU6502.scala 19:21 66:22]
  wire  _GEN_928 = 8'h86 == opcode ? flagN : _GEN_910; // @[CPU6502.scala 31:22 66:22]
  wire  _GEN_929 = 8'h86 == opcode ? flagZ : _GEN_911; // @[CPU6502.scala 26:22 66:22]
  wire [7:0] _GEN_930 = 8'h86 == opcode ? regSP : _GEN_912; // @[CPU6502.scala 21:22 66:22]
  wire [7:0] _GEN_931 = 8'h86 == opcode ? regA : _GEN_913; // @[CPU6502.scala 18:21 66:22]
  wire  _GEN_932 = 8'h86 == opcode ? flagC : _GEN_914; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_933 = 8'h86 == opcode ? flagI : _GEN_915; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_934 = 8'h86 == opcode ? flagD : _GEN_916; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_935 = 8'h86 == opcode ? flagV : _GEN_917; // @[CPU6502.scala 30:22 66:22]
  wire [15:0] _GEN_937 = 8'hc6 == opcode ? _GEN_204 : _GEN_919; // @[CPU6502.scala 66:22]
  wire  _GEN_938 = 8'hc6 == opcode ? _GEN_14 : _GEN_920; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_939 = 8'hc6 == opcode ? _GEN_15 : _GEN_921; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_940 = 8'hc6 == opcode ? _GEN_5 : _GEN_922; // @[CPU6502.scala 66:22]
  wire [2:0] _GEN_941 = 8'hc6 == opcode ? _GEN_208 : _GEN_923; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_942 = 8'hc6 == opcode ? _GEN_339 : _GEN_924; // @[CPU6502.scala 66:22]
  wire  _GEN_943 = 8'hc6 == opcode ? _GEN_211 : _GEN_925; // @[CPU6502.scala 66:22]
  wire  _GEN_944 = 8'hc6 == opcode ? _GEN_341 : _GEN_928; // @[CPU6502.scala 66:22]
  wire  _GEN_945 = 8'hc6 == opcode ? _GEN_342 : _GEN_929; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_946 = 8'hc6 == opcode ? _GEN_214 : _GEN_926; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_947 = 8'hc6 == opcode ? regX : _GEN_927; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_948 = 8'hc6 == opcode ? regSP : _GEN_930; // @[CPU6502.scala 21:22 66:22]
  wire [7:0] _GEN_949 = 8'hc6 == opcode ? regA : _GEN_931; // @[CPU6502.scala 18:21 66:22]
  wire  _GEN_950 = 8'hc6 == opcode ? flagC : _GEN_932; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_951 = 8'hc6 == opcode ? flagI : _GEN_933; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_952 = 8'hc6 == opcode ? flagD : _GEN_934; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_953 = 8'hc6 == opcode ? flagV : _GEN_935; // @[CPU6502.scala 30:22 66:22]
  wire [15:0] _GEN_955 = 8'he6 == opcode ? _GEN_204 : _GEN_937; // @[CPU6502.scala 66:22]
  wire  _GEN_956 = 8'he6 == opcode ? _GEN_14 : _GEN_938; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_957 = 8'he6 == opcode ? _GEN_15 : _GEN_939; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_958 = 8'he6 == opcode ? _GEN_5 : _GEN_940; // @[CPU6502.scala 66:22]
  wire [2:0] _GEN_959 = 8'he6 == opcode ? _GEN_208 : _GEN_941; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_960 = 8'he6 == opcode ? _GEN_315 : _GEN_942; // @[CPU6502.scala 66:22]
  wire  _GEN_961 = 8'he6 == opcode ? _GEN_211 : _GEN_943; // @[CPU6502.scala 66:22]
  wire  _GEN_962 = 8'he6 == opcode ? _GEN_317 : _GEN_944; // @[CPU6502.scala 66:22]
  wire  _GEN_963 = 8'he6 == opcode ? _GEN_318 : _GEN_945; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_964 = 8'he6 == opcode ? _GEN_214 : _GEN_946; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_965 = 8'he6 == opcode ? regX : _GEN_947; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_966 = 8'he6 == opcode ? regSP : _GEN_948; // @[CPU6502.scala 21:22 66:22]
  wire [7:0] _GEN_967 = 8'he6 == opcode ? regA : _GEN_949; // @[CPU6502.scala 18:21 66:22]
  wire  _GEN_968 = 8'he6 == opcode ? flagC : _GEN_950; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_969 = 8'he6 == opcode ? flagI : _GEN_951; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_970 = 8'he6 == opcode ? flagD : _GEN_952; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_971 = 8'he6 == opcode ? flagV : _GEN_953; // @[CPU6502.scala 30:22 66:22]
  wire [15:0] _GEN_973 = 8'h66 == opcode ? _GEN_204 : _GEN_955; // @[CPU6502.scala 66:22]
  wire  _GEN_974 = 8'h66 == opcode ? _GEN_14 : _GEN_956; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_975 = 8'h66 == opcode ? _GEN_15 : _GEN_957; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_976 = 8'h66 == opcode ? _GEN_5 : _GEN_958; // @[CPU6502.scala 66:22]
  wire [2:0] _GEN_977 = 8'h66 == opcode ? _GEN_208 : _GEN_959; // @[CPU6502.scala 66:22]
  wire  _GEN_978 = 8'h66 == opcode ? _GEN_236 : _GEN_968; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_979 = 8'h66 == opcode ? _GEN_291 : _GEN_960; // @[CPU6502.scala 66:22]
  wire  _GEN_980 = 8'h66 == opcode ? _GEN_211 : _GEN_961; // @[CPU6502.scala 66:22]
  wire  _GEN_981 = 8'h66 == opcode ? _GEN_293 : _GEN_962; // @[CPU6502.scala 66:22]
  wire  _GEN_982 = 8'h66 == opcode ? _GEN_294 : _GEN_963; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_983 = 8'h66 == opcode ? _GEN_214 : _GEN_964; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_984 = 8'h66 == opcode ? regX : _GEN_965; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_985 = 8'h66 == opcode ? regSP : _GEN_966; // @[CPU6502.scala 21:22 66:22]
  wire [7:0] _GEN_986 = 8'h66 == opcode ? regA : _GEN_967; // @[CPU6502.scala 18:21 66:22]
  wire  _GEN_987 = 8'h66 == opcode ? flagI : _GEN_969; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_988 = 8'h66 == opcode ? flagD : _GEN_970; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_989 = 8'h66 == opcode ? flagV : _GEN_971; // @[CPU6502.scala 30:22 66:22]
  wire  _GEN_991 = 8'h6a == opcode ? regA[0] : _GEN_978; // @[CPU6502.scala 627:17 66:22]
  wire [7:0] _GEN_992 = 8'h6a == opcode ? result_17 : _GEN_986; // @[CPU6502.scala 629:16 66:22]
  wire  _GEN_993 = 8'h6a == opcode ? result_17[7] : _GEN_981; // @[CPU6502.scala 50:11 66:22]
  wire  _GEN_994 = 8'h6a == opcode ? result_17 == 8'h0 : _GEN_982; // @[CPU6502.scala 51:11 66:22]
  wire [1:0] _GEN_995 = 8'h6a == opcode ? 2'h0 : _GEN_983; // @[CPU6502.scala 631:17 66:22]
  wire [15:0] _GEN_996 = 8'h6a == opcode ? regPC : _GEN_973; // @[CPU6502.scala 42:14 66:22]
  wire  _GEN_997 = 8'h6a == opcode ? 1'h0 : _GEN_974; // @[CPU6502.scala 45:14 66:22]
  wire [15:0] _GEN_998 = 8'h6a == opcode ? operand : _GEN_975; // @[CPU6502.scala 66:22 38:24]
  wire [15:0] _GEN_999 = 8'h6a == opcode ? regPC : _GEN_976; // @[CPU6502.scala 22:22 66:22]
  wire [2:0] _GEN_1000 = 8'h6a == opcode ? cycle : _GEN_977; // @[CPU6502.scala 39:22 66:22]
  wire [7:0] _GEN_1001 = 8'h6a == opcode ? 8'h0 : _GEN_979; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1002 = 8'h6a == opcode ? 1'h0 : _GEN_980; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_1003 = 8'h6a == opcode ? regX : _GEN_984; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_1004 = 8'h6a == opcode ? regSP : _GEN_985; // @[CPU6502.scala 21:22 66:22]
  wire  _GEN_1005 = 8'h6a == opcode ? flagI : _GEN_987; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_1006 = 8'h6a == opcode ? flagD : _GEN_988; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_1007 = 8'h6a == opcode ? flagV : _GEN_989; // @[CPU6502.scala 30:22 66:22]
  wire [15:0] _GEN_1009 = 8'h26 == opcode ? _GEN_204 : _GEN_996; // @[CPU6502.scala 66:22]
  wire  _GEN_1010 = 8'h26 == opcode ? _GEN_14 : _GEN_997; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_1011 = 8'h26 == opcode ? _GEN_15 : _GEN_998; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_1012 = 8'h26 == opcode ? _GEN_5 : _GEN_999; // @[CPU6502.scala 66:22]
  wire [2:0] _GEN_1013 = 8'h26 == opcode ? _GEN_208 : _GEN_1000; // @[CPU6502.scala 66:22]
  wire  _GEN_1014 = 8'h26 == opcode ? _GEN_209 : _GEN_991; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_1015 = 8'h26 == opcode ? _GEN_264 : _GEN_1001; // @[CPU6502.scala 66:22]
  wire  _GEN_1016 = 8'h26 == opcode ? _GEN_211 : _GEN_1002; // @[CPU6502.scala 66:22]
  wire  _GEN_1017 = 8'h26 == opcode ? _GEN_266 : _GEN_993; // @[CPU6502.scala 66:22]
  wire  _GEN_1018 = 8'h26 == opcode ? _GEN_267 : _GEN_994; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_1019 = 8'h26 == opcode ? _GEN_214 : _GEN_995; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_1020 = 8'h26 == opcode ? regA : _GEN_992; // @[CPU6502.scala 18:21 66:22]
  wire [7:0] _GEN_1021 = 8'h26 == opcode ? regX : _GEN_1003; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_1022 = 8'h26 == opcode ? regSP : _GEN_1004; // @[CPU6502.scala 21:22 66:22]
  wire  _GEN_1023 = 8'h26 == opcode ? flagI : _GEN_1005; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_1024 = 8'h26 == opcode ? flagD : _GEN_1006; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_1025 = 8'h26 == opcode ? flagV : _GEN_1007; // @[CPU6502.scala 30:22 66:22]
  wire  _GEN_1027 = 8'h2a == opcode ? regA[7] : _GEN_1014; // @[CPU6502.scala 592:17 66:22]
  wire [7:0] _GEN_1028 = 8'h2a == opcode ? result_15 : _GEN_1020; // @[CPU6502.scala 594:16 66:22]
  wire  _GEN_1029 = 8'h2a == opcode ? result_15[7] : _GEN_1017; // @[CPU6502.scala 50:11 66:22]
  wire  _GEN_1030 = 8'h2a == opcode ? result_15 == 8'h0 : _GEN_1018; // @[CPU6502.scala 51:11 66:22]
  wire [1:0] _GEN_1031 = 8'h2a == opcode ? 2'h0 : _GEN_1019; // @[CPU6502.scala 596:17 66:22]
  wire [15:0] _GEN_1032 = 8'h2a == opcode ? regPC : _GEN_1009; // @[CPU6502.scala 42:14 66:22]
  wire  _GEN_1033 = 8'h2a == opcode ? 1'h0 : _GEN_1010; // @[CPU6502.scala 45:14 66:22]
  wire [15:0] _GEN_1034 = 8'h2a == opcode ? operand : _GEN_1011; // @[CPU6502.scala 66:22 38:24]
  wire [15:0] _GEN_1035 = 8'h2a == opcode ? regPC : _GEN_1012; // @[CPU6502.scala 22:22 66:22]
  wire [2:0] _GEN_1036 = 8'h2a == opcode ? cycle : _GEN_1013; // @[CPU6502.scala 39:22 66:22]
  wire [7:0] _GEN_1037 = 8'h2a == opcode ? 8'h0 : _GEN_1015; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1038 = 8'h2a == opcode ? 1'h0 : _GEN_1016; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_1039 = 8'h2a == opcode ? regX : _GEN_1021; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_1040 = 8'h2a == opcode ? regSP : _GEN_1022; // @[CPU6502.scala 21:22 66:22]
  wire  _GEN_1041 = 8'h2a == opcode ? flagI : _GEN_1023; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_1042 = 8'h2a == opcode ? flagD : _GEN_1024; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_1043 = 8'h2a == opcode ? flagV : _GEN_1025; // @[CPU6502.scala 30:22 66:22]
  wire [15:0] _GEN_1045 = 8'h46 == opcode ? _GEN_204 : _GEN_1032; // @[CPU6502.scala 66:22]
  wire  _GEN_1046 = 8'h46 == opcode ? _GEN_14 : _GEN_1033; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_1047 = 8'h46 == opcode ? _GEN_15 : _GEN_1034; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_1048 = 8'h46 == opcode ? _GEN_5 : _GEN_1035; // @[CPU6502.scala 66:22]
  wire [2:0] _GEN_1049 = 8'h46 == opcode ? _GEN_208 : _GEN_1036; // @[CPU6502.scala 66:22]
  wire  _GEN_1050 = 8'h46 == opcode ? _GEN_236 : _GEN_1027; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_1051 = 8'h46 == opcode ? _GEN_237 : _GEN_1037; // @[CPU6502.scala 66:22]
  wire  _GEN_1052 = 8'h46 == opcode ? _GEN_211 : _GEN_1038; // @[CPU6502.scala 66:22]
  wire  _GEN_1053 = 8'h46 == opcode ? _GEN_239 : _GEN_1029; // @[CPU6502.scala 66:22]
  wire  _GEN_1054 = 8'h46 == opcode ? _GEN_240 : _GEN_1030; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_1055 = 8'h46 == opcode ? _GEN_214 : _GEN_1031; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_1056 = 8'h46 == opcode ? regA : _GEN_1028; // @[CPU6502.scala 18:21 66:22]
  wire [7:0] _GEN_1057 = 8'h46 == opcode ? regX : _GEN_1039; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_1058 = 8'h46 == opcode ? regSP : _GEN_1040; // @[CPU6502.scala 21:22 66:22]
  wire  _GEN_1059 = 8'h46 == opcode ? flagI : _GEN_1041; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_1060 = 8'h46 == opcode ? flagD : _GEN_1042; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_1061 = 8'h46 == opcode ? flagV : _GEN_1043; // @[CPU6502.scala 30:22 66:22]
  wire  _GEN_1063 = 8'h4a == opcode ? regA[0] : _GEN_1050; // @[CPU6502.scala 558:17 66:22]
  wire [7:0] _GEN_1064 = 8'h4a == opcode ? result_13 : _GEN_1056; // @[CPU6502.scala 560:16 66:22]
  wire  _GEN_1065 = 8'h4a == opcode ? result_13[7] : _GEN_1053; // @[CPU6502.scala 50:11 66:22]
  wire  _GEN_1066 = 8'h4a == opcode ? result_13 == 8'h0 : _GEN_1054; // @[CPU6502.scala 51:11 66:22]
  wire [1:0] _GEN_1067 = 8'h4a == opcode ? 2'h0 : _GEN_1055; // @[CPU6502.scala 562:17 66:22]
  wire [15:0] _GEN_1068 = 8'h4a == opcode ? regPC : _GEN_1045; // @[CPU6502.scala 42:14 66:22]
  wire  _GEN_1069 = 8'h4a == opcode ? 1'h0 : _GEN_1046; // @[CPU6502.scala 45:14 66:22]
  wire [15:0] _GEN_1070 = 8'h4a == opcode ? operand : _GEN_1047; // @[CPU6502.scala 66:22 38:24]
  wire [15:0] _GEN_1071 = 8'h4a == opcode ? regPC : _GEN_1048; // @[CPU6502.scala 22:22 66:22]
  wire [2:0] _GEN_1072 = 8'h4a == opcode ? cycle : _GEN_1049; // @[CPU6502.scala 39:22 66:22]
  wire [7:0] _GEN_1073 = 8'h4a == opcode ? 8'h0 : _GEN_1051; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1074 = 8'h4a == opcode ? 1'h0 : _GEN_1052; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_1075 = 8'h4a == opcode ? regX : _GEN_1057; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_1076 = 8'h4a == opcode ? regSP : _GEN_1058; // @[CPU6502.scala 21:22 66:22]
  wire  _GEN_1077 = 8'h4a == opcode ? flagI : _GEN_1059; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_1078 = 8'h4a == opcode ? flagD : _GEN_1060; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_1079 = 8'h4a == opcode ? flagV : _GEN_1061; // @[CPU6502.scala 30:22 66:22]
  wire [15:0] _GEN_1081 = 8'h6 == opcode ? _GEN_204 : _GEN_1068; // @[CPU6502.scala 66:22]
  wire  _GEN_1082 = 8'h6 == opcode ? _GEN_14 : _GEN_1069; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_1083 = 8'h6 == opcode ? _GEN_15 : _GEN_1070; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_1084 = 8'h6 == opcode ? _GEN_5 : _GEN_1071; // @[CPU6502.scala 66:22]
  wire [2:0] _GEN_1085 = 8'h6 == opcode ? _GEN_208 : _GEN_1072; // @[CPU6502.scala 66:22]
  wire  _GEN_1086 = 8'h6 == opcode ? _GEN_209 : _GEN_1063; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_1087 = 8'h6 == opcode ? _GEN_210 : _GEN_1073; // @[CPU6502.scala 66:22]
  wire  _GEN_1088 = 8'h6 == opcode ? _GEN_211 : _GEN_1074; // @[CPU6502.scala 66:22]
  wire  _GEN_1089 = 8'h6 == opcode ? _GEN_212 : _GEN_1065; // @[CPU6502.scala 66:22]
  wire  _GEN_1090 = 8'h6 == opcode ? _GEN_213 : _GEN_1066; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_1091 = 8'h6 == opcode ? _GEN_214 : _GEN_1067; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_1092 = 8'h6 == opcode ? regA : _GEN_1064; // @[CPU6502.scala 18:21 66:22]
  wire [7:0] _GEN_1093 = 8'h6 == opcode ? regX : _GEN_1075; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_1094 = 8'h6 == opcode ? regSP : _GEN_1076; // @[CPU6502.scala 21:22 66:22]
  wire  _GEN_1095 = 8'h6 == opcode ? flagI : _GEN_1077; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_1096 = 8'h6 == opcode ? flagD : _GEN_1078; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_1097 = 8'h6 == opcode ? flagV : _GEN_1079; // @[CPU6502.scala 30:22 66:22]
  wire  _GEN_1099 = 8'ha == opcode ? regA[7] : _GEN_1086; // @[CPU6502.scala 524:17 66:22]
  wire [7:0] _GEN_1100 = 8'ha == opcode ? result_11 : _GEN_1092; // @[CPU6502.scala 527:16 66:22]
  wire  _GEN_1101 = 8'ha == opcode ? result_11[7] : _GEN_1089; // @[CPU6502.scala 50:11 66:22]
  wire  _GEN_1102 = 8'ha == opcode ? result_11 == 8'h0 : _GEN_1090; // @[CPU6502.scala 51:11 66:22]
  wire [1:0] _GEN_1103 = 8'ha == opcode ? 2'h0 : _GEN_1091; // @[CPU6502.scala 529:17 66:22]
  wire [15:0] _GEN_1104 = 8'ha == opcode ? regPC : _GEN_1081; // @[CPU6502.scala 42:14 66:22]
  wire  _GEN_1105 = 8'ha == opcode ? 1'h0 : _GEN_1082; // @[CPU6502.scala 45:14 66:22]
  wire [15:0] _GEN_1106 = 8'ha == opcode ? operand : _GEN_1083; // @[CPU6502.scala 66:22 38:24]
  wire [15:0] _GEN_1107 = 8'ha == opcode ? regPC : _GEN_1084; // @[CPU6502.scala 22:22 66:22]
  wire [2:0] _GEN_1108 = 8'ha == opcode ? cycle : _GEN_1085; // @[CPU6502.scala 39:22 66:22]
  wire [7:0] _GEN_1109 = 8'ha == opcode ? 8'h0 : _GEN_1087; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1110 = 8'ha == opcode ? 1'h0 : _GEN_1088; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_1111 = 8'ha == opcode ? regX : _GEN_1093; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_1112 = 8'ha == opcode ? regSP : _GEN_1094; // @[CPU6502.scala 21:22 66:22]
  wire  _GEN_1113 = 8'ha == opcode ? flagI : _GEN_1095; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_1114 = 8'ha == opcode ? flagD : _GEN_1096; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_1115 = 8'ha == opcode ? flagV : _GEN_1097; // @[CPU6502.scala 30:22 66:22]
  wire [15:0] _GEN_1117 = 8'h24 == opcode ? _GEN_13 : _GEN_1104; // @[CPU6502.scala 66:22]
  wire  _GEN_1118 = 8'h24 == opcode ? _GEN_14 : _GEN_1105; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_1119 = 8'h24 == opcode ? _GEN_15 : _GEN_1106; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_1120 = 8'h24 == opcode ? _GEN_5 : _GEN_1107; // @[CPU6502.scala 66:22]
  wire [2:0] _GEN_1121 = 8'h24 == opcode ? _GEN_17 : _GEN_1108; // @[CPU6502.scala 66:22]
  wire  _GEN_1122 = 8'h24 == opcode ? _GEN_184 : _GEN_1102; // @[CPU6502.scala 66:22]
  wire  _GEN_1123 = 8'h24 == opcode ? _GEN_19 : _GEN_1101; // @[CPU6502.scala 66:22]
  wire  _GEN_1124 = 8'h24 == opcode ? _GEN_186 : _GEN_1115; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_1125 = 8'h24 == opcode ? _GEN_21 : _GEN_1103; // @[CPU6502.scala 66:22]
  wire  _GEN_1126 = 8'h24 == opcode ? flagC : _GEN_1099; // @[CPU6502.scala 25:22 66:22]
  wire [7:0] _GEN_1127 = 8'h24 == opcode ? regA : _GEN_1100; // @[CPU6502.scala 18:21 66:22]
  wire [7:0] _GEN_1128 = 8'h24 == opcode ? 8'h0 : _GEN_1109; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1129 = 8'h24 == opcode ? 1'h0 : _GEN_1110; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_1130 = 8'h24 == opcode ? regX : _GEN_1111; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_1131 = 8'h24 == opcode ? regSP : _GEN_1112; // @[CPU6502.scala 21:22 66:22]
  wire  _GEN_1132 = 8'h24 == opcode ? flagI : _GEN_1113; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_1133 = 8'h24 == opcode ? flagD : _GEN_1114; // @[CPU6502.scala 28:22 66:22]
  wire [15:0] _GEN_1135 = 8'hc0 == opcode ? regPC : _GEN_1117; // @[CPU6502.scala 66:22]
  wire  _GEN_1136 = 8'hc0 == opcode ? _T_3 : _GEN_1118; // @[CPU6502.scala 66:22]
  wire  _GEN_1137 = 8'hc0 == opcode ? _GEN_168 : _GEN_1126; // @[CPU6502.scala 66:22]
  wire  _GEN_1138 = 8'hc0 == opcode ? _GEN_169 : _GEN_1122; // @[CPU6502.scala 66:22]
  wire  _GEN_1139 = 8'hc0 == opcode ? _GEN_170 : _GEN_1123; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_1140 = 8'hc0 == opcode ? _GEN_5 : _GEN_1120; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_1141 = 8'hc0 == opcode ? _GEN_6 : _GEN_1125; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_1142 = 8'hc0 == opcode ? operand : _GEN_1119; // @[CPU6502.scala 66:22 38:24]
  wire [2:0] _GEN_1143 = 8'hc0 == opcode ? cycle : _GEN_1121; // @[CPU6502.scala 39:22 66:22]
  wire  _GEN_1144 = 8'hc0 == opcode ? flagV : _GEN_1124; // @[CPU6502.scala 30:22 66:22]
  wire [7:0] _GEN_1145 = 8'hc0 == opcode ? regA : _GEN_1127; // @[CPU6502.scala 18:21 66:22]
  wire [7:0] _GEN_1146 = 8'hc0 == opcode ? 8'h0 : _GEN_1128; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1147 = 8'hc0 == opcode ? 1'h0 : _GEN_1129; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_1148 = 8'hc0 == opcode ? regX : _GEN_1130; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_1149 = 8'hc0 == opcode ? regSP : _GEN_1131; // @[CPU6502.scala 21:22 66:22]
  wire  _GEN_1150 = 8'hc0 == opcode ? flagI : _GEN_1132; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_1151 = 8'hc0 == opcode ? flagD : _GEN_1133; // @[CPU6502.scala 28:22 66:22]
  wire [15:0] _GEN_1153 = 8'he0 == opcode ? regPC : _GEN_1135; // @[CPU6502.scala 66:22]
  wire  _GEN_1154 = 8'he0 == opcode ? _T_3 : _GEN_1136; // @[CPU6502.scala 66:22]
  wire  _GEN_1155 = 8'he0 == opcode ? _GEN_161 : _GEN_1137; // @[CPU6502.scala 66:22]
  wire  _GEN_1156 = 8'he0 == opcode ? _GEN_162 : _GEN_1138; // @[CPU6502.scala 66:22]
  wire  _GEN_1157 = 8'he0 == opcode ? _GEN_163 : _GEN_1139; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_1158 = 8'he0 == opcode ? _GEN_5 : _GEN_1140; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_1159 = 8'he0 == opcode ? _GEN_6 : _GEN_1141; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_1160 = 8'he0 == opcode ? operand : _GEN_1142; // @[CPU6502.scala 66:22 38:24]
  wire [2:0] _GEN_1161 = 8'he0 == opcode ? cycle : _GEN_1143; // @[CPU6502.scala 39:22 66:22]
  wire  _GEN_1162 = 8'he0 == opcode ? flagV : _GEN_1144; // @[CPU6502.scala 30:22 66:22]
  wire [7:0] _GEN_1163 = 8'he0 == opcode ? regA : _GEN_1145; // @[CPU6502.scala 18:21 66:22]
  wire [7:0] _GEN_1164 = 8'he0 == opcode ? 8'h0 : _GEN_1146; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1165 = 8'he0 == opcode ? 1'h0 : _GEN_1147; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_1166 = 8'he0 == opcode ? regX : _GEN_1148; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_1167 = 8'he0 == opcode ? regSP : _GEN_1149; // @[CPU6502.scala 21:22 66:22]
  wire  _GEN_1168 = 8'he0 == opcode ? flagI : _GEN_1150; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_1169 = 8'he0 == opcode ? flagD : _GEN_1151; // @[CPU6502.scala 28:22 66:22]
  wire [15:0] _GEN_1171 = 8'hc5 == opcode ? _GEN_13 : _GEN_1153; // @[CPU6502.scala 66:22]
  wire  _GEN_1172 = 8'hc5 == opcode ? _GEN_14 : _GEN_1154; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_1173 = 8'hc5 == opcode ? _GEN_15 : _GEN_1160; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_1174 = 8'hc5 == opcode ? _GEN_5 : _GEN_1158; // @[CPU6502.scala 66:22]
  wire [2:0] _GEN_1175 = 8'hc5 == opcode ? _GEN_17 : _GEN_1161; // @[CPU6502.scala 66:22]
  wire  _GEN_1176 = 8'hc5 == opcode ? _GEN_155 : _GEN_1155; // @[CPU6502.scala 66:22]
  wire  _GEN_1177 = 8'hc5 == opcode ? _GEN_156 : _GEN_1156; // @[CPU6502.scala 66:22]
  wire  _GEN_1178 = 8'hc5 == opcode ? _GEN_157 : _GEN_1157; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_1179 = 8'hc5 == opcode ? _GEN_21 : _GEN_1159; // @[CPU6502.scala 66:22]
  wire  _GEN_1180 = 8'hc5 == opcode ? flagV : _GEN_1162; // @[CPU6502.scala 30:22 66:22]
  wire [7:0] _GEN_1181 = 8'hc5 == opcode ? regA : _GEN_1163; // @[CPU6502.scala 18:21 66:22]
  wire [7:0] _GEN_1182 = 8'hc5 == opcode ? 8'h0 : _GEN_1164; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1183 = 8'hc5 == opcode ? 1'h0 : _GEN_1165; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_1184 = 8'hc5 == opcode ? regX : _GEN_1166; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_1185 = 8'hc5 == opcode ? regSP : _GEN_1167; // @[CPU6502.scala 21:22 66:22]
  wire  _GEN_1186 = 8'hc5 == opcode ? flagI : _GEN_1168; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_1187 = 8'hc5 == opcode ? flagD : _GEN_1169; // @[CPU6502.scala 28:22 66:22]
  wire [15:0] _GEN_1189 = 8'hc9 == opcode ? regPC : _GEN_1171; // @[CPU6502.scala 66:22]
  wire  _GEN_1190 = 8'hc9 == opcode ? _T_3 : _GEN_1172; // @[CPU6502.scala 66:22]
  wire  _GEN_1191 = 8'hc9 == opcode ? _GEN_139 : _GEN_1176; // @[CPU6502.scala 66:22]
  wire  _GEN_1192 = 8'hc9 == opcode ? _GEN_140 : _GEN_1177; // @[CPU6502.scala 66:22]
  wire  _GEN_1193 = 8'hc9 == opcode ? _GEN_141 : _GEN_1178; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_1194 = 8'hc9 == opcode ? _GEN_5 : _GEN_1174; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_1195 = 8'hc9 == opcode ? _GEN_6 : _GEN_1179; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_1196 = 8'hc9 == opcode ? operand : _GEN_1173; // @[CPU6502.scala 66:22 38:24]
  wire [2:0] _GEN_1197 = 8'hc9 == opcode ? cycle : _GEN_1175; // @[CPU6502.scala 39:22 66:22]
  wire  _GEN_1198 = 8'hc9 == opcode ? flagV : _GEN_1180; // @[CPU6502.scala 30:22 66:22]
  wire [7:0] _GEN_1199 = 8'hc9 == opcode ? regA : _GEN_1181; // @[CPU6502.scala 18:21 66:22]
  wire [7:0] _GEN_1200 = 8'hc9 == opcode ? 8'h0 : _GEN_1182; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1201 = 8'hc9 == opcode ? 1'h0 : _GEN_1183; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_1202 = 8'hc9 == opcode ? regX : _GEN_1184; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_1203 = 8'hc9 == opcode ? regSP : _GEN_1185; // @[CPU6502.scala 21:22 66:22]
  wire  _GEN_1204 = 8'hc9 == opcode ? flagI : _GEN_1186; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_1205 = 8'hc9 == opcode ? flagD : _GEN_1187; // @[CPU6502.scala 28:22 66:22]
  wire [15:0] _GEN_1207 = 8'h70 == opcode ? regPC : _GEN_1189; // @[CPU6502.scala 66:22]
  wire  _GEN_1208 = 8'h70 == opcode ? _T_3 : _GEN_1190; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_1209 = 8'h70 == opcode ? _GEN_135 : _GEN_1194; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_1210 = 8'h70 == opcode ? _GEN_6 : _GEN_1195; // @[CPU6502.scala 66:22]
  wire  _GEN_1211 = 8'h70 == opcode ? flagC : _GEN_1191; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_1212 = 8'h70 == opcode ? flagZ : _GEN_1192; // @[CPU6502.scala 26:22 66:22]
  wire  _GEN_1213 = 8'h70 == opcode ? flagN : _GEN_1193; // @[CPU6502.scala 31:22 66:22]
  wire [15:0] _GEN_1214 = 8'h70 == opcode ? operand : _GEN_1196; // @[CPU6502.scala 66:22 38:24]
  wire [2:0] _GEN_1215 = 8'h70 == opcode ? cycle : _GEN_1197; // @[CPU6502.scala 39:22 66:22]
  wire  _GEN_1216 = 8'h70 == opcode ? flagV : _GEN_1198; // @[CPU6502.scala 30:22 66:22]
  wire [7:0] _GEN_1217 = 8'h70 == opcode ? regA : _GEN_1199; // @[CPU6502.scala 18:21 66:22]
  wire [7:0] _GEN_1218 = 8'h70 == opcode ? 8'h0 : _GEN_1200; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1219 = 8'h70 == opcode ? 1'h0 : _GEN_1201; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_1220 = 8'h70 == opcode ? regX : _GEN_1202; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_1221 = 8'h70 == opcode ? regSP : _GEN_1203; // @[CPU6502.scala 21:22 66:22]
  wire  _GEN_1222 = 8'h70 == opcode ? flagI : _GEN_1204; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_1223 = 8'h70 == opcode ? flagD : _GEN_1205; // @[CPU6502.scala 28:22 66:22]
  wire [15:0] _GEN_1225 = 8'h50 == opcode ? regPC : _GEN_1207; // @[CPU6502.scala 66:22]
  wire  _GEN_1226 = 8'h50 == opcode ? _T_3 : _GEN_1208; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_1227 = 8'h50 == opcode ? _GEN_130 : _GEN_1209; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_1228 = 8'h50 == opcode ? _GEN_6 : _GEN_1210; // @[CPU6502.scala 66:22]
  wire  _GEN_1229 = 8'h50 == opcode ? flagC : _GEN_1211; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_1230 = 8'h50 == opcode ? flagZ : _GEN_1212; // @[CPU6502.scala 26:22 66:22]
  wire  _GEN_1231 = 8'h50 == opcode ? flagN : _GEN_1213; // @[CPU6502.scala 31:22 66:22]
  wire [15:0] _GEN_1232 = 8'h50 == opcode ? operand : _GEN_1214; // @[CPU6502.scala 66:22 38:24]
  wire [2:0] _GEN_1233 = 8'h50 == opcode ? cycle : _GEN_1215; // @[CPU6502.scala 39:22 66:22]
  wire  _GEN_1234 = 8'h50 == opcode ? flagV : _GEN_1216; // @[CPU6502.scala 30:22 66:22]
  wire [7:0] _GEN_1235 = 8'h50 == opcode ? regA : _GEN_1217; // @[CPU6502.scala 18:21 66:22]
  wire [7:0] _GEN_1236 = 8'h50 == opcode ? 8'h0 : _GEN_1218; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1237 = 8'h50 == opcode ? 1'h0 : _GEN_1219; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_1238 = 8'h50 == opcode ? regX : _GEN_1220; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_1239 = 8'h50 == opcode ? regSP : _GEN_1221; // @[CPU6502.scala 21:22 66:22]
  wire  _GEN_1240 = 8'h50 == opcode ? flagI : _GEN_1222; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_1241 = 8'h50 == opcode ? flagD : _GEN_1223; // @[CPU6502.scala 28:22 66:22]
  wire [15:0] _GEN_1243 = 8'h10 == opcode ? regPC : _GEN_1225; // @[CPU6502.scala 66:22]
  wire  _GEN_1244 = 8'h10 == opcode ? _T_3 : _GEN_1226; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_1245 = 8'h10 == opcode ? _GEN_125 : _GEN_1227; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_1246 = 8'h10 == opcode ? _GEN_6 : _GEN_1228; // @[CPU6502.scala 66:22]
  wire  _GEN_1247 = 8'h10 == opcode ? flagC : _GEN_1229; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_1248 = 8'h10 == opcode ? flagZ : _GEN_1230; // @[CPU6502.scala 26:22 66:22]
  wire  _GEN_1249 = 8'h10 == opcode ? flagN : _GEN_1231; // @[CPU6502.scala 31:22 66:22]
  wire [15:0] _GEN_1250 = 8'h10 == opcode ? operand : _GEN_1232; // @[CPU6502.scala 66:22 38:24]
  wire [2:0] _GEN_1251 = 8'h10 == opcode ? cycle : _GEN_1233; // @[CPU6502.scala 39:22 66:22]
  wire  _GEN_1252 = 8'h10 == opcode ? flagV : _GEN_1234; // @[CPU6502.scala 30:22 66:22]
  wire [7:0] _GEN_1253 = 8'h10 == opcode ? regA : _GEN_1235; // @[CPU6502.scala 18:21 66:22]
  wire [7:0] _GEN_1254 = 8'h10 == opcode ? 8'h0 : _GEN_1236; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1255 = 8'h10 == opcode ? 1'h0 : _GEN_1237; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_1256 = 8'h10 == opcode ? regX : _GEN_1238; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_1257 = 8'h10 == opcode ? regSP : _GEN_1239; // @[CPU6502.scala 21:22 66:22]
  wire  _GEN_1258 = 8'h10 == opcode ? flagI : _GEN_1240; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_1259 = 8'h10 == opcode ? flagD : _GEN_1241; // @[CPU6502.scala 28:22 66:22]
  wire [15:0] _GEN_1261 = 8'h30 == opcode ? regPC : _GEN_1243; // @[CPU6502.scala 66:22]
  wire  _GEN_1262 = 8'h30 == opcode ? _T_3 : _GEN_1244; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_1263 = 8'h30 == opcode ? _GEN_120 : _GEN_1245; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_1264 = 8'h30 == opcode ? _GEN_6 : _GEN_1246; // @[CPU6502.scala 66:22]
  wire  _GEN_1265 = 8'h30 == opcode ? flagC : _GEN_1247; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_1266 = 8'h30 == opcode ? flagZ : _GEN_1248; // @[CPU6502.scala 26:22 66:22]
  wire  _GEN_1267 = 8'h30 == opcode ? flagN : _GEN_1249; // @[CPU6502.scala 31:22 66:22]
  wire [15:0] _GEN_1268 = 8'h30 == opcode ? operand : _GEN_1250; // @[CPU6502.scala 66:22 38:24]
  wire [2:0] _GEN_1269 = 8'h30 == opcode ? cycle : _GEN_1251; // @[CPU6502.scala 39:22 66:22]
  wire  _GEN_1270 = 8'h30 == opcode ? flagV : _GEN_1252; // @[CPU6502.scala 30:22 66:22]
  wire [7:0] _GEN_1271 = 8'h30 == opcode ? regA : _GEN_1253; // @[CPU6502.scala 18:21 66:22]
  wire [7:0] _GEN_1272 = 8'h30 == opcode ? 8'h0 : _GEN_1254; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1273 = 8'h30 == opcode ? 1'h0 : _GEN_1255; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_1274 = 8'h30 == opcode ? regX : _GEN_1256; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_1275 = 8'h30 == opcode ? regSP : _GEN_1257; // @[CPU6502.scala 21:22 66:22]
  wire  _GEN_1276 = 8'h30 == opcode ? flagI : _GEN_1258; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_1277 = 8'h30 == opcode ? flagD : _GEN_1259; // @[CPU6502.scala 28:22 66:22]
  wire [15:0] _GEN_1279 = 8'h90 == opcode ? regPC : _GEN_1261; // @[CPU6502.scala 66:22]
  wire  _GEN_1280 = 8'h90 == opcode ? _T_3 : _GEN_1262; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_1281 = 8'h90 == opcode ? _GEN_115 : _GEN_1263; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_1282 = 8'h90 == opcode ? _GEN_6 : _GEN_1264; // @[CPU6502.scala 66:22]
  wire  _GEN_1283 = 8'h90 == opcode ? flagC : _GEN_1265; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_1284 = 8'h90 == opcode ? flagZ : _GEN_1266; // @[CPU6502.scala 26:22 66:22]
  wire  _GEN_1285 = 8'h90 == opcode ? flagN : _GEN_1267; // @[CPU6502.scala 31:22 66:22]
  wire [15:0] _GEN_1286 = 8'h90 == opcode ? operand : _GEN_1268; // @[CPU6502.scala 66:22 38:24]
  wire [2:0] _GEN_1287 = 8'h90 == opcode ? cycle : _GEN_1269; // @[CPU6502.scala 39:22 66:22]
  wire  _GEN_1288 = 8'h90 == opcode ? flagV : _GEN_1270; // @[CPU6502.scala 30:22 66:22]
  wire [7:0] _GEN_1289 = 8'h90 == opcode ? regA : _GEN_1271; // @[CPU6502.scala 18:21 66:22]
  wire [7:0] _GEN_1290 = 8'h90 == opcode ? 8'h0 : _GEN_1272; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1291 = 8'h90 == opcode ? 1'h0 : _GEN_1273; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_1292 = 8'h90 == opcode ? regX : _GEN_1274; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_1293 = 8'h90 == opcode ? regSP : _GEN_1275; // @[CPU6502.scala 21:22 66:22]
  wire  _GEN_1294 = 8'h90 == opcode ? flagI : _GEN_1276; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_1295 = 8'h90 == opcode ? flagD : _GEN_1277; // @[CPU6502.scala 28:22 66:22]
  wire [15:0] _GEN_1297 = 8'hb0 == opcode ? regPC : _GEN_1279; // @[CPU6502.scala 66:22]
  wire  _GEN_1298 = 8'hb0 == opcode ? _T_3 : _GEN_1280; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_1299 = 8'hb0 == opcode ? _GEN_110 : _GEN_1281; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_1300 = 8'hb0 == opcode ? _GEN_6 : _GEN_1282; // @[CPU6502.scala 66:22]
  wire  _GEN_1301 = 8'hb0 == opcode ? flagC : _GEN_1283; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_1302 = 8'hb0 == opcode ? flagZ : _GEN_1284; // @[CPU6502.scala 26:22 66:22]
  wire  _GEN_1303 = 8'hb0 == opcode ? flagN : _GEN_1285; // @[CPU6502.scala 31:22 66:22]
  wire [15:0] _GEN_1304 = 8'hb0 == opcode ? operand : _GEN_1286; // @[CPU6502.scala 66:22 38:24]
  wire [2:0] _GEN_1305 = 8'hb0 == opcode ? cycle : _GEN_1287; // @[CPU6502.scala 39:22 66:22]
  wire  _GEN_1306 = 8'hb0 == opcode ? flagV : _GEN_1288; // @[CPU6502.scala 30:22 66:22]
  wire [7:0] _GEN_1307 = 8'hb0 == opcode ? regA : _GEN_1289; // @[CPU6502.scala 18:21 66:22]
  wire [7:0] _GEN_1308 = 8'hb0 == opcode ? 8'h0 : _GEN_1290; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1309 = 8'hb0 == opcode ? 1'h0 : _GEN_1291; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_1310 = 8'hb0 == opcode ? regX : _GEN_1292; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_1311 = 8'hb0 == opcode ? regSP : _GEN_1293; // @[CPU6502.scala 21:22 66:22]
  wire  _GEN_1312 = 8'hb0 == opcode ? flagI : _GEN_1294; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_1313 = 8'hb0 == opcode ? flagD : _GEN_1295; // @[CPU6502.scala 28:22 66:22]
  wire [15:0] _GEN_1315 = 8'hd0 == opcode ? regPC : _GEN_1297; // @[CPU6502.scala 66:22]
  wire  _GEN_1316 = 8'hd0 == opcode ? _T_3 : _GEN_1298; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_1317 = 8'hd0 == opcode ? _GEN_105 : _GEN_1299; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_1318 = 8'hd0 == opcode ? _GEN_6 : _GEN_1300; // @[CPU6502.scala 66:22]
  wire  _GEN_1319 = 8'hd0 == opcode ? flagC : _GEN_1301; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_1320 = 8'hd0 == opcode ? flagZ : _GEN_1302; // @[CPU6502.scala 26:22 66:22]
  wire  _GEN_1321 = 8'hd0 == opcode ? flagN : _GEN_1303; // @[CPU6502.scala 31:22 66:22]
  wire [15:0] _GEN_1322 = 8'hd0 == opcode ? operand : _GEN_1304; // @[CPU6502.scala 66:22 38:24]
  wire [2:0] _GEN_1323 = 8'hd0 == opcode ? cycle : _GEN_1305; // @[CPU6502.scala 39:22 66:22]
  wire  _GEN_1324 = 8'hd0 == opcode ? flagV : _GEN_1306; // @[CPU6502.scala 30:22 66:22]
  wire [7:0] _GEN_1325 = 8'hd0 == opcode ? regA : _GEN_1307; // @[CPU6502.scala 18:21 66:22]
  wire [7:0] _GEN_1326 = 8'hd0 == opcode ? 8'h0 : _GEN_1308; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1327 = 8'hd0 == opcode ? 1'h0 : _GEN_1309; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_1328 = 8'hd0 == opcode ? regX : _GEN_1310; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_1329 = 8'hd0 == opcode ? regSP : _GEN_1311; // @[CPU6502.scala 21:22 66:22]
  wire  _GEN_1330 = 8'hd0 == opcode ? flagI : _GEN_1312; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_1331 = 8'hd0 == opcode ? flagD : _GEN_1313; // @[CPU6502.scala 28:22 66:22]
  wire [15:0] _GEN_1333 = 8'hf0 == opcode ? regPC : _GEN_1315; // @[CPU6502.scala 66:22]
  wire  _GEN_1334 = 8'hf0 == opcode ? _T_3 : _GEN_1316; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_1335 = 8'hf0 == opcode ? _GEN_100 : _GEN_1317; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_1336 = 8'hf0 == opcode ? _GEN_6 : _GEN_1318; // @[CPU6502.scala 66:22]
  wire  _GEN_1337 = 8'hf0 == opcode ? flagC : _GEN_1319; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_1338 = 8'hf0 == opcode ? flagZ : _GEN_1320; // @[CPU6502.scala 26:22 66:22]
  wire  _GEN_1339 = 8'hf0 == opcode ? flagN : _GEN_1321; // @[CPU6502.scala 31:22 66:22]
  wire [15:0] _GEN_1340 = 8'hf0 == opcode ? operand : _GEN_1322; // @[CPU6502.scala 66:22 38:24]
  wire [2:0] _GEN_1341 = 8'hf0 == opcode ? cycle : _GEN_1323; // @[CPU6502.scala 39:22 66:22]
  wire  _GEN_1342 = 8'hf0 == opcode ? flagV : _GEN_1324; // @[CPU6502.scala 30:22 66:22]
  wire [7:0] _GEN_1343 = 8'hf0 == opcode ? regA : _GEN_1325; // @[CPU6502.scala 18:21 66:22]
  wire [7:0] _GEN_1344 = 8'hf0 == opcode ? 8'h0 : _GEN_1326; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1345 = 8'hf0 == opcode ? 1'h0 : _GEN_1327; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_1346 = 8'hf0 == opcode ? regX : _GEN_1328; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_1347 = 8'hf0 == opcode ? regSP : _GEN_1329; // @[CPU6502.scala 21:22 66:22]
  wire  _GEN_1348 = 8'hf0 == opcode ? flagI : _GEN_1330; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_1349 = 8'hf0 == opcode ? flagD : _GEN_1331; // @[CPU6502.scala 28:22 66:22]
  wire [15:0] _GEN_1351 = 8'h4c == opcode ? regPC : _GEN_1333; // @[CPU6502.scala 66:22]
  wire  _GEN_1352 = 8'h4c == opcode ? _GEN_14 : _GEN_1334; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_1353 = 8'h4c == opcode ? _GEN_15 : _GEN_1340; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_1354 = 8'h4c == opcode ? _GEN_94 : _GEN_1335; // @[CPU6502.scala 66:22]
  wire [2:0] _GEN_1355 = 8'h4c == opcode ? _GEN_17 : _GEN_1341; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_1356 = 8'h4c == opcode ? _GEN_21 : _GEN_1336; // @[CPU6502.scala 66:22]
  wire  _GEN_1357 = 8'h4c == opcode ? flagC : _GEN_1337; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_1358 = 8'h4c == opcode ? flagZ : _GEN_1338; // @[CPU6502.scala 26:22 66:22]
  wire  _GEN_1359 = 8'h4c == opcode ? flagN : _GEN_1339; // @[CPU6502.scala 31:22 66:22]
  wire  _GEN_1360 = 8'h4c == opcode ? flagV : _GEN_1342; // @[CPU6502.scala 30:22 66:22]
  wire [7:0] _GEN_1361 = 8'h4c == opcode ? regA : _GEN_1343; // @[CPU6502.scala 18:21 66:22]
  wire [7:0] _GEN_1362 = 8'h4c == opcode ? 8'h0 : _GEN_1344; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1363 = 8'h4c == opcode ? 1'h0 : _GEN_1345; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_1364 = 8'h4c == opcode ? regX : _GEN_1346; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_1365 = 8'h4c == opcode ? regSP : _GEN_1347; // @[CPU6502.scala 21:22 66:22]
  wire  _GEN_1366 = 8'h4c == opcode ? flagI : _GEN_1348; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_1367 = 8'h4c == opcode ? flagD : _GEN_1349; // @[CPU6502.scala 28:22 66:22]
  wire [1:0] _GEN_1369 = 8'hea == opcode ? 2'h0 : _GEN_1356; // @[CPU6502.scala 311:17 66:22]
  wire [15:0] _GEN_1370 = 8'hea == opcode ? regPC : _GEN_1351; // @[CPU6502.scala 42:14 66:22]
  wire  _GEN_1371 = 8'hea == opcode ? 1'h0 : _GEN_1352; // @[CPU6502.scala 45:14 66:22]
  wire [15:0] _GEN_1372 = 8'hea == opcode ? operand : _GEN_1353; // @[CPU6502.scala 66:22 38:24]
  wire [15:0] _GEN_1373 = 8'hea == opcode ? regPC : _GEN_1354; // @[CPU6502.scala 22:22 66:22]
  wire [2:0] _GEN_1374 = 8'hea == opcode ? cycle : _GEN_1355; // @[CPU6502.scala 39:22 66:22]
  wire  _GEN_1375 = 8'hea == opcode ? flagC : _GEN_1357; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_1376 = 8'hea == opcode ? flagZ : _GEN_1358; // @[CPU6502.scala 26:22 66:22]
  wire  _GEN_1377 = 8'hea == opcode ? flagN : _GEN_1359; // @[CPU6502.scala 31:22 66:22]
  wire  _GEN_1378 = 8'hea == opcode ? flagV : _GEN_1360; // @[CPU6502.scala 30:22 66:22]
  wire [7:0] _GEN_1379 = 8'hea == opcode ? regA : _GEN_1361; // @[CPU6502.scala 18:21 66:22]
  wire [7:0] _GEN_1380 = 8'hea == opcode ? 8'h0 : _GEN_1362; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1381 = 8'hea == opcode ? 1'h0 : _GEN_1363; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_1382 = 8'hea == opcode ? regX : _GEN_1364; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_1383 = 8'hea == opcode ? regSP : _GEN_1365; // @[CPU6502.scala 21:22 66:22]
  wire  _GEN_1384 = 8'hea == opcode ? flagI : _GEN_1366; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_1385 = 8'hea == opcode ? flagD : _GEN_1367; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_1387 = 8'hb8 == opcode ? 1'h0 : _GEN_1378; // @[CPU6502.scala 305:17 66:22]
  wire [1:0] _GEN_1388 = 8'hb8 == opcode ? 2'h0 : _GEN_1369; // @[CPU6502.scala 306:17 66:22]
  wire [15:0] _GEN_1389 = 8'hb8 == opcode ? regPC : _GEN_1370; // @[CPU6502.scala 42:14 66:22]
  wire  _GEN_1390 = 8'hb8 == opcode ? 1'h0 : _GEN_1371; // @[CPU6502.scala 45:14 66:22]
  wire [15:0] _GEN_1391 = 8'hb8 == opcode ? operand : _GEN_1372; // @[CPU6502.scala 66:22 38:24]
  wire [15:0] _GEN_1392 = 8'hb8 == opcode ? regPC : _GEN_1373; // @[CPU6502.scala 22:22 66:22]
  wire [2:0] _GEN_1393 = 8'hb8 == opcode ? cycle : _GEN_1374; // @[CPU6502.scala 39:22 66:22]
  wire  _GEN_1394 = 8'hb8 == opcode ? flagC : _GEN_1375; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_1395 = 8'hb8 == opcode ? flagZ : _GEN_1376; // @[CPU6502.scala 26:22 66:22]
  wire  _GEN_1396 = 8'hb8 == opcode ? flagN : _GEN_1377; // @[CPU6502.scala 31:22 66:22]
  wire [7:0] _GEN_1397 = 8'hb8 == opcode ? regA : _GEN_1379; // @[CPU6502.scala 18:21 66:22]
  wire [7:0] _GEN_1398 = 8'hb8 == opcode ? 8'h0 : _GEN_1380; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1399 = 8'hb8 == opcode ? 1'h0 : _GEN_1381; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_1400 = 8'hb8 == opcode ? regX : _GEN_1382; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_1401 = 8'hb8 == opcode ? regSP : _GEN_1383; // @[CPU6502.scala 21:22 66:22]
  wire  _GEN_1402 = 8'hb8 == opcode ? flagI : _GEN_1384; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_1403 = 8'hb8 == opcode ? flagD : _GEN_1385; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_1405 = 8'h78 == opcode | _GEN_1402; // @[CPU6502.scala 299:17 66:22]
  wire [1:0] _GEN_1406 = 8'h78 == opcode ? 2'h0 : _GEN_1388; // @[CPU6502.scala 300:17 66:22]
  wire  _GEN_1407 = 8'h78 == opcode ? flagV : _GEN_1387; // @[CPU6502.scala 30:22 66:22]
  wire [15:0] _GEN_1408 = 8'h78 == opcode ? regPC : _GEN_1389; // @[CPU6502.scala 42:14 66:22]
  wire  _GEN_1409 = 8'h78 == opcode ? 1'h0 : _GEN_1390; // @[CPU6502.scala 45:14 66:22]
  wire [15:0] _GEN_1410 = 8'h78 == opcode ? operand : _GEN_1391; // @[CPU6502.scala 66:22 38:24]
  wire [15:0] _GEN_1411 = 8'h78 == opcode ? regPC : _GEN_1392; // @[CPU6502.scala 22:22 66:22]
  wire [2:0] _GEN_1412 = 8'h78 == opcode ? cycle : _GEN_1393; // @[CPU6502.scala 39:22 66:22]
  wire  _GEN_1413 = 8'h78 == opcode ? flagC : _GEN_1394; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_1414 = 8'h78 == opcode ? flagZ : _GEN_1395; // @[CPU6502.scala 26:22 66:22]
  wire  _GEN_1415 = 8'h78 == opcode ? flagN : _GEN_1396; // @[CPU6502.scala 31:22 66:22]
  wire [7:0] _GEN_1416 = 8'h78 == opcode ? regA : _GEN_1397; // @[CPU6502.scala 18:21 66:22]
  wire [7:0] _GEN_1417 = 8'h78 == opcode ? 8'h0 : _GEN_1398; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1418 = 8'h78 == opcode ? 1'h0 : _GEN_1399; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_1419 = 8'h78 == opcode ? regX : _GEN_1400; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_1420 = 8'h78 == opcode ? regSP : _GEN_1401; // @[CPU6502.scala 21:22 66:22]
  wire  _GEN_1421 = 8'h78 == opcode ? flagD : _GEN_1403; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_1423 = 8'h58 == opcode ? 1'h0 : _GEN_1405; // @[CPU6502.scala 293:17 66:22]
  wire [1:0] _GEN_1424 = 8'h58 == opcode ? 2'h0 : _GEN_1406; // @[CPU6502.scala 294:17 66:22]
  wire  _GEN_1425 = 8'h58 == opcode ? flagV : _GEN_1407; // @[CPU6502.scala 30:22 66:22]
  wire [15:0] _GEN_1426 = 8'h58 == opcode ? regPC : _GEN_1408; // @[CPU6502.scala 42:14 66:22]
  wire  _GEN_1427 = 8'h58 == opcode ? 1'h0 : _GEN_1409; // @[CPU6502.scala 45:14 66:22]
  wire [15:0] _GEN_1428 = 8'h58 == opcode ? operand : _GEN_1410; // @[CPU6502.scala 66:22 38:24]
  wire [15:0] _GEN_1429 = 8'h58 == opcode ? regPC : _GEN_1411; // @[CPU6502.scala 22:22 66:22]
  wire [2:0] _GEN_1430 = 8'h58 == opcode ? cycle : _GEN_1412; // @[CPU6502.scala 39:22 66:22]
  wire  _GEN_1431 = 8'h58 == opcode ? flagC : _GEN_1413; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_1432 = 8'h58 == opcode ? flagZ : _GEN_1414; // @[CPU6502.scala 26:22 66:22]
  wire  _GEN_1433 = 8'h58 == opcode ? flagN : _GEN_1415; // @[CPU6502.scala 31:22 66:22]
  wire [7:0] _GEN_1434 = 8'h58 == opcode ? regA : _GEN_1416; // @[CPU6502.scala 18:21 66:22]
  wire [7:0] _GEN_1435 = 8'h58 == opcode ? 8'h0 : _GEN_1417; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1436 = 8'h58 == opcode ? 1'h0 : _GEN_1418; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_1437 = 8'h58 == opcode ? regX : _GEN_1419; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_1438 = 8'h58 == opcode ? regSP : _GEN_1420; // @[CPU6502.scala 21:22 66:22]
  wire  _GEN_1439 = 8'h58 == opcode ? flagD : _GEN_1421; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_1441 = 8'hf8 == opcode | _GEN_1439; // @[CPU6502.scala 287:17 66:22]
  wire [1:0] _GEN_1442 = 8'hf8 == opcode ? 2'h0 : _GEN_1424; // @[CPU6502.scala 288:17 66:22]
  wire  _GEN_1443 = 8'hf8 == opcode ? flagI : _GEN_1423; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_1444 = 8'hf8 == opcode ? flagV : _GEN_1425; // @[CPU6502.scala 30:22 66:22]
  wire [15:0] _GEN_1445 = 8'hf8 == opcode ? regPC : _GEN_1426; // @[CPU6502.scala 42:14 66:22]
  wire  _GEN_1446 = 8'hf8 == opcode ? 1'h0 : _GEN_1427; // @[CPU6502.scala 45:14 66:22]
  wire [15:0] _GEN_1447 = 8'hf8 == opcode ? operand : _GEN_1428; // @[CPU6502.scala 66:22 38:24]
  wire [15:0] _GEN_1448 = 8'hf8 == opcode ? regPC : _GEN_1429; // @[CPU6502.scala 22:22 66:22]
  wire [2:0] _GEN_1449 = 8'hf8 == opcode ? cycle : _GEN_1430; // @[CPU6502.scala 39:22 66:22]
  wire  _GEN_1450 = 8'hf8 == opcode ? flagC : _GEN_1431; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_1451 = 8'hf8 == opcode ? flagZ : _GEN_1432; // @[CPU6502.scala 26:22 66:22]
  wire  _GEN_1452 = 8'hf8 == opcode ? flagN : _GEN_1433; // @[CPU6502.scala 31:22 66:22]
  wire [7:0] _GEN_1453 = 8'hf8 == opcode ? regA : _GEN_1434; // @[CPU6502.scala 18:21 66:22]
  wire [7:0] _GEN_1454 = 8'hf8 == opcode ? 8'h0 : _GEN_1435; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1455 = 8'hf8 == opcode ? 1'h0 : _GEN_1436; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_1456 = 8'hf8 == opcode ? regX : _GEN_1437; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_1457 = 8'hf8 == opcode ? regSP : _GEN_1438; // @[CPU6502.scala 21:22 66:22]
  wire  _GEN_1459 = 8'hd8 == opcode ? 1'h0 : _GEN_1441; // @[CPU6502.scala 281:17 66:22]
  wire [1:0] _GEN_1460 = 8'hd8 == opcode ? 2'h0 : _GEN_1442; // @[CPU6502.scala 282:17 66:22]
  wire  _GEN_1461 = 8'hd8 == opcode ? flagI : _GEN_1443; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_1462 = 8'hd8 == opcode ? flagV : _GEN_1444; // @[CPU6502.scala 30:22 66:22]
  wire [15:0] _GEN_1463 = 8'hd8 == opcode ? regPC : _GEN_1445; // @[CPU6502.scala 42:14 66:22]
  wire  _GEN_1464 = 8'hd8 == opcode ? 1'h0 : _GEN_1446; // @[CPU6502.scala 45:14 66:22]
  wire [15:0] _GEN_1465 = 8'hd8 == opcode ? operand : _GEN_1447; // @[CPU6502.scala 66:22 38:24]
  wire [15:0] _GEN_1466 = 8'hd8 == opcode ? regPC : _GEN_1448; // @[CPU6502.scala 22:22 66:22]
  wire [2:0] _GEN_1467 = 8'hd8 == opcode ? cycle : _GEN_1449; // @[CPU6502.scala 39:22 66:22]
  wire  _GEN_1468 = 8'hd8 == opcode ? flagC : _GEN_1450; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_1469 = 8'hd8 == opcode ? flagZ : _GEN_1451; // @[CPU6502.scala 26:22 66:22]
  wire  _GEN_1470 = 8'hd8 == opcode ? flagN : _GEN_1452; // @[CPU6502.scala 31:22 66:22]
  wire [7:0] _GEN_1471 = 8'hd8 == opcode ? regA : _GEN_1453; // @[CPU6502.scala 18:21 66:22]
  wire [7:0] _GEN_1472 = 8'hd8 == opcode ? 8'h0 : _GEN_1454; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1473 = 8'hd8 == opcode ? 1'h0 : _GEN_1455; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_1474 = 8'hd8 == opcode ? regX : _GEN_1456; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_1475 = 8'hd8 == opcode ? regSP : _GEN_1457; // @[CPU6502.scala 21:22 66:22]
  wire  _GEN_1477 = 8'h38 == opcode | _GEN_1468; // @[CPU6502.scala 275:17 66:22]
  wire [1:0] _GEN_1478 = 8'h38 == opcode ? 2'h0 : _GEN_1460; // @[CPU6502.scala 276:17 66:22]
  wire  _GEN_1479 = 8'h38 == opcode ? flagD : _GEN_1459; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_1480 = 8'h38 == opcode ? flagI : _GEN_1461; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_1481 = 8'h38 == opcode ? flagV : _GEN_1462; // @[CPU6502.scala 30:22 66:22]
  wire [15:0] _GEN_1482 = 8'h38 == opcode ? regPC : _GEN_1463; // @[CPU6502.scala 42:14 66:22]
  wire  _GEN_1483 = 8'h38 == opcode ? 1'h0 : _GEN_1464; // @[CPU6502.scala 45:14 66:22]
  wire [15:0] _GEN_1484 = 8'h38 == opcode ? operand : _GEN_1465; // @[CPU6502.scala 66:22 38:24]
  wire [15:0] _GEN_1485 = 8'h38 == opcode ? regPC : _GEN_1466; // @[CPU6502.scala 22:22 66:22]
  wire [2:0] _GEN_1486 = 8'h38 == opcode ? cycle : _GEN_1467; // @[CPU6502.scala 39:22 66:22]
  wire  _GEN_1487 = 8'h38 == opcode ? flagZ : _GEN_1469; // @[CPU6502.scala 26:22 66:22]
  wire  _GEN_1488 = 8'h38 == opcode ? flagN : _GEN_1470; // @[CPU6502.scala 31:22 66:22]
  wire [7:0] _GEN_1489 = 8'h38 == opcode ? regA : _GEN_1471; // @[CPU6502.scala 18:21 66:22]
  wire [7:0] _GEN_1490 = 8'h38 == opcode ? 8'h0 : _GEN_1472; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1491 = 8'h38 == opcode ? 1'h0 : _GEN_1473; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_1492 = 8'h38 == opcode ? regX : _GEN_1474; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_1493 = 8'h38 == opcode ? regSP : _GEN_1475; // @[CPU6502.scala 21:22 66:22]
  wire  _GEN_1495 = 8'h18 == opcode ? 1'h0 : _GEN_1477; // @[CPU6502.scala 269:17 66:22]
  wire [1:0] _GEN_1496 = 8'h18 == opcode ? 2'h0 : _GEN_1478; // @[CPU6502.scala 270:17 66:22]
  wire  _GEN_1497 = 8'h18 == opcode ? flagD : _GEN_1479; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_1498 = 8'h18 == opcode ? flagI : _GEN_1480; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_1499 = 8'h18 == opcode ? flagV : _GEN_1481; // @[CPU6502.scala 30:22 66:22]
  wire [15:0] _GEN_1500 = 8'h18 == opcode ? regPC : _GEN_1482; // @[CPU6502.scala 42:14 66:22]
  wire  _GEN_1501 = 8'h18 == opcode ? 1'h0 : _GEN_1483; // @[CPU6502.scala 45:14 66:22]
  wire [15:0] _GEN_1502 = 8'h18 == opcode ? operand : _GEN_1484; // @[CPU6502.scala 66:22 38:24]
  wire [15:0] _GEN_1503 = 8'h18 == opcode ? regPC : _GEN_1485; // @[CPU6502.scala 22:22 66:22]
  wire [2:0] _GEN_1504 = 8'h18 == opcode ? cycle : _GEN_1486; // @[CPU6502.scala 39:22 66:22]
  wire  _GEN_1505 = 8'h18 == opcode ? flagZ : _GEN_1487; // @[CPU6502.scala 26:22 66:22]
  wire  _GEN_1506 = 8'h18 == opcode ? flagN : _GEN_1488; // @[CPU6502.scala 31:22 66:22]
  wire [7:0] _GEN_1507 = 8'h18 == opcode ? regA : _GEN_1489; // @[CPU6502.scala 18:21 66:22]
  wire [7:0] _GEN_1508 = 8'h18 == opcode ? 8'h0 : _GEN_1490; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1509 = 8'h18 == opcode ? 1'h0 : _GEN_1491; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_1510 = 8'h18 == opcode ? regX : _GEN_1492; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_1511 = 8'h18 == opcode ? regSP : _GEN_1493; // @[CPU6502.scala 21:22 66:22]
  wire [7:0] _GEN_1513 = 8'h98 == opcode ? regY : _GEN_1507; // @[CPU6502.scala 262:16 66:22]
  wire  _GEN_1514 = 8'h98 == opcode ? regY[7] : _GEN_1506; // @[CPU6502.scala 50:11 66:22]
  wire  _GEN_1515 = 8'h98 == opcode ? regY == 8'h0 : _GEN_1505; // @[CPU6502.scala 51:11 66:22]
  wire [1:0] _GEN_1516 = 8'h98 == opcode ? 2'h0 : _GEN_1496; // @[CPU6502.scala 264:17 66:22]
  wire  _GEN_1517 = 8'h98 == opcode ? flagC : _GEN_1495; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_1518 = 8'h98 == opcode ? flagD : _GEN_1497; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_1519 = 8'h98 == opcode ? flagI : _GEN_1498; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_1520 = 8'h98 == opcode ? flagV : _GEN_1499; // @[CPU6502.scala 30:22 66:22]
  wire [15:0] _GEN_1521 = 8'h98 == opcode ? regPC : _GEN_1500; // @[CPU6502.scala 42:14 66:22]
  wire  _GEN_1522 = 8'h98 == opcode ? 1'h0 : _GEN_1501; // @[CPU6502.scala 45:14 66:22]
  wire [15:0] _GEN_1523 = 8'h98 == opcode ? operand : _GEN_1502; // @[CPU6502.scala 66:22 38:24]
  wire [15:0] _GEN_1524 = 8'h98 == opcode ? regPC : _GEN_1503; // @[CPU6502.scala 22:22 66:22]
  wire [2:0] _GEN_1525 = 8'h98 == opcode ? cycle : _GEN_1504; // @[CPU6502.scala 39:22 66:22]
  wire [7:0] _GEN_1526 = 8'h98 == opcode ? 8'h0 : _GEN_1508; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1527 = 8'h98 == opcode ? 1'h0 : _GEN_1509; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_1528 = 8'h98 == opcode ? regX : _GEN_1510; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_1529 = 8'h98 == opcode ? regSP : _GEN_1511; // @[CPU6502.scala 21:22 66:22]
  wire [7:0] _GEN_1531 = 8'h8a == opcode ? regX : _GEN_1513; // @[CPU6502.scala 255:16 66:22]
  wire  _GEN_1532 = 8'h8a == opcode ? regX[7] : _GEN_1514; // @[CPU6502.scala 50:11 66:22]
  wire  _GEN_1533 = 8'h8a == opcode ? regX == 8'h0 : _GEN_1515; // @[CPU6502.scala 51:11 66:22]
  wire [1:0] _GEN_1534 = 8'h8a == opcode ? 2'h0 : _GEN_1516; // @[CPU6502.scala 257:17 66:22]
  wire  _GEN_1535 = 8'h8a == opcode ? flagC : _GEN_1517; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_1536 = 8'h8a == opcode ? flagD : _GEN_1518; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_1537 = 8'h8a == opcode ? flagI : _GEN_1519; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_1538 = 8'h8a == opcode ? flagV : _GEN_1520; // @[CPU6502.scala 30:22 66:22]
  wire [15:0] _GEN_1539 = 8'h8a == opcode ? regPC : _GEN_1521; // @[CPU6502.scala 42:14 66:22]
  wire  _GEN_1540 = 8'h8a == opcode ? 1'h0 : _GEN_1522; // @[CPU6502.scala 45:14 66:22]
  wire [15:0] _GEN_1541 = 8'h8a == opcode ? operand : _GEN_1523; // @[CPU6502.scala 66:22 38:24]
  wire [15:0] _GEN_1542 = 8'h8a == opcode ? regPC : _GEN_1524; // @[CPU6502.scala 22:22 66:22]
  wire [2:0] _GEN_1543 = 8'h8a == opcode ? cycle : _GEN_1525; // @[CPU6502.scala 39:22 66:22]
  wire [7:0] _GEN_1544 = 8'h8a == opcode ? 8'h0 : _GEN_1526; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1545 = 8'h8a == opcode ? 1'h0 : _GEN_1527; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_1546 = 8'h8a == opcode ? regX : _GEN_1528; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_1547 = 8'h8a == opcode ? regSP : _GEN_1529; // @[CPU6502.scala 21:22 66:22]
  wire [7:0] _GEN_1549 = 8'ha8 == opcode ? regA : regY; // @[CPU6502.scala 248:16 20:21 66:22]
  wire  _GEN_1550 = 8'ha8 == opcode ? regA[7] : _GEN_1532; // @[CPU6502.scala 50:11 66:22]
  wire  _GEN_1551 = 8'ha8 == opcode ? regA == 8'h0 : _GEN_1533; // @[CPU6502.scala 51:11 66:22]
  wire [1:0] _GEN_1552 = 8'ha8 == opcode ? 2'h0 : _GEN_1534; // @[CPU6502.scala 250:17 66:22]
  wire [7:0] _GEN_1553 = 8'ha8 == opcode ? regA : _GEN_1531; // @[CPU6502.scala 18:21 66:22]
  wire  _GEN_1554 = 8'ha8 == opcode ? flagC : _GEN_1535; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_1555 = 8'ha8 == opcode ? flagD : _GEN_1536; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_1556 = 8'ha8 == opcode ? flagI : _GEN_1537; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_1557 = 8'ha8 == opcode ? flagV : _GEN_1538; // @[CPU6502.scala 30:22 66:22]
  wire [15:0] _GEN_1558 = 8'ha8 == opcode ? regPC : _GEN_1539; // @[CPU6502.scala 42:14 66:22]
  wire  _GEN_1559 = 8'ha8 == opcode ? 1'h0 : _GEN_1540; // @[CPU6502.scala 45:14 66:22]
  wire [15:0] _GEN_1560 = 8'ha8 == opcode ? operand : _GEN_1541; // @[CPU6502.scala 66:22 38:24]
  wire [15:0] _GEN_1561 = 8'ha8 == opcode ? regPC : _GEN_1542; // @[CPU6502.scala 22:22 66:22]
  wire [2:0] _GEN_1562 = 8'ha8 == opcode ? cycle : _GEN_1543; // @[CPU6502.scala 39:22 66:22]
  wire [7:0] _GEN_1563 = 8'ha8 == opcode ? 8'h0 : _GEN_1544; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1564 = 8'ha8 == opcode ? 1'h0 : _GEN_1545; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_1565 = 8'ha8 == opcode ? regX : _GEN_1546; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_1566 = 8'ha8 == opcode ? regSP : _GEN_1547; // @[CPU6502.scala 21:22 66:22]
  wire [7:0] _GEN_1568 = 8'haa == opcode ? regA : _GEN_1565; // @[CPU6502.scala 241:16 66:22]
  wire  _GEN_1569 = 8'haa == opcode ? regA[7] : _GEN_1550; // @[CPU6502.scala 50:11 66:22]
  wire  _GEN_1570 = 8'haa == opcode ? regA == 8'h0 : _GEN_1551; // @[CPU6502.scala 51:11 66:22]
  wire [1:0] _GEN_1571 = 8'haa == opcode ? 2'h0 : _GEN_1552; // @[CPU6502.scala 243:17 66:22]
  wire [7:0] _GEN_1572 = 8'haa == opcode ? regY : _GEN_1549; // @[CPU6502.scala 20:21 66:22]
  wire [7:0] _GEN_1573 = 8'haa == opcode ? regA : _GEN_1553; // @[CPU6502.scala 18:21 66:22]
  wire  _GEN_1574 = 8'haa == opcode ? flagC : _GEN_1554; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_1575 = 8'haa == opcode ? flagD : _GEN_1555; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_1576 = 8'haa == opcode ? flagI : _GEN_1556; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_1577 = 8'haa == opcode ? flagV : _GEN_1557; // @[CPU6502.scala 30:22 66:22]
  wire [15:0] _GEN_1578 = 8'haa == opcode ? regPC : _GEN_1558; // @[CPU6502.scala 42:14 66:22]
  wire  _GEN_1579 = 8'haa == opcode ? 1'h0 : _GEN_1559; // @[CPU6502.scala 45:14 66:22]
  wire [15:0] _GEN_1580 = 8'haa == opcode ? operand : _GEN_1560; // @[CPU6502.scala 66:22 38:24]
  wire [15:0] _GEN_1581 = 8'haa == opcode ? regPC : _GEN_1561; // @[CPU6502.scala 22:22 66:22]
  wire [2:0] _GEN_1582 = 8'haa == opcode ? cycle : _GEN_1562; // @[CPU6502.scala 39:22 66:22]
  wire [7:0] _GEN_1583 = 8'haa == opcode ? 8'h0 : _GEN_1563; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1584 = 8'haa == opcode ? 1'h0 : _GEN_1564; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_1585 = 8'haa == opcode ? regSP : _GEN_1566; // @[CPU6502.scala 21:22 66:22]
  wire [7:0] _GEN_1587 = 8'h88 == opcode ? result_6 : _GEN_1572; // @[CPU6502.scala 234:16 66:22]
  wire  _GEN_1588 = 8'h88 == opcode ? result_6[7] : _GEN_1569; // @[CPU6502.scala 50:11 66:22]
  wire  _GEN_1589 = 8'h88 == opcode ? result_6 == 8'h0 : _GEN_1570; // @[CPU6502.scala 51:11 66:22]
  wire [1:0] _GEN_1590 = 8'h88 == opcode ? 2'h0 : _GEN_1571; // @[CPU6502.scala 236:17 66:22]
  wire [7:0] _GEN_1591 = 8'h88 == opcode ? regX : _GEN_1568; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_1592 = 8'h88 == opcode ? regA : _GEN_1573; // @[CPU6502.scala 18:21 66:22]
  wire  _GEN_1593 = 8'h88 == opcode ? flagC : _GEN_1574; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_1594 = 8'h88 == opcode ? flagD : _GEN_1575; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_1595 = 8'h88 == opcode ? flagI : _GEN_1576; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_1596 = 8'h88 == opcode ? flagV : _GEN_1577; // @[CPU6502.scala 30:22 66:22]
  wire [15:0] _GEN_1597 = 8'h88 == opcode ? regPC : _GEN_1578; // @[CPU6502.scala 42:14 66:22]
  wire  _GEN_1598 = 8'h88 == opcode ? 1'h0 : _GEN_1579; // @[CPU6502.scala 45:14 66:22]
  wire [15:0] _GEN_1599 = 8'h88 == opcode ? operand : _GEN_1580; // @[CPU6502.scala 66:22 38:24]
  wire [15:0] _GEN_1600 = 8'h88 == opcode ? regPC : _GEN_1581; // @[CPU6502.scala 22:22 66:22]
  wire [2:0] _GEN_1601 = 8'h88 == opcode ? cycle : _GEN_1582; // @[CPU6502.scala 39:22 66:22]
  wire [7:0] _GEN_1602 = 8'h88 == opcode ? 8'h0 : _GEN_1583; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1603 = 8'h88 == opcode ? 1'h0 : _GEN_1584; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_1604 = 8'h88 == opcode ? regSP : _GEN_1585; // @[CPU6502.scala 21:22 66:22]
  wire [7:0] _GEN_1606 = 8'hca == opcode ? result_5 : _GEN_1591; // @[CPU6502.scala 226:16 66:22]
  wire  _GEN_1607 = 8'hca == opcode ? result_5[7] : _GEN_1588; // @[CPU6502.scala 50:11 66:22]
  wire  _GEN_1608 = 8'hca == opcode ? result_5 == 8'h0 : _GEN_1589; // @[CPU6502.scala 51:11 66:22]
  wire [1:0] _GEN_1609 = 8'hca == opcode ? 2'h0 : _GEN_1590; // @[CPU6502.scala 228:17 66:22]
  wire [7:0] _GEN_1610 = 8'hca == opcode ? regY : _GEN_1587; // @[CPU6502.scala 20:21 66:22]
  wire [7:0] _GEN_1611 = 8'hca == opcode ? regA : _GEN_1592; // @[CPU6502.scala 18:21 66:22]
  wire  _GEN_1612 = 8'hca == opcode ? flagC : _GEN_1593; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_1613 = 8'hca == opcode ? flagD : _GEN_1594; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_1614 = 8'hca == opcode ? flagI : _GEN_1595; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_1615 = 8'hca == opcode ? flagV : _GEN_1596; // @[CPU6502.scala 30:22 66:22]
  wire [15:0] _GEN_1616 = 8'hca == opcode ? regPC : _GEN_1597; // @[CPU6502.scala 42:14 66:22]
  wire  _GEN_1617 = 8'hca == opcode ? 1'h0 : _GEN_1598; // @[CPU6502.scala 45:14 66:22]
  wire [15:0] _GEN_1618 = 8'hca == opcode ? operand : _GEN_1599; // @[CPU6502.scala 66:22 38:24]
  wire [15:0] _GEN_1619 = 8'hca == opcode ? regPC : _GEN_1600; // @[CPU6502.scala 22:22 66:22]
  wire [2:0] _GEN_1620 = 8'hca == opcode ? cycle : _GEN_1601; // @[CPU6502.scala 39:22 66:22]
  wire [7:0] _GEN_1621 = 8'hca == opcode ? 8'h0 : _GEN_1602; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1622 = 8'hca == opcode ? 1'h0 : _GEN_1603; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_1623 = 8'hca == opcode ? regSP : _GEN_1604; // @[CPU6502.scala 21:22 66:22]
  wire [7:0] _GEN_1625 = 8'hc8 == opcode ? result_4 : _GEN_1610; // @[CPU6502.scala 218:16 66:22]
  wire  _GEN_1626 = 8'hc8 == opcode ? result_4[7] : _GEN_1607; // @[CPU6502.scala 50:11 66:22]
  wire  _GEN_1627 = 8'hc8 == opcode ? result_4 == 8'h0 : _GEN_1608; // @[CPU6502.scala 51:11 66:22]
  wire [1:0] _GEN_1628 = 8'hc8 == opcode ? 2'h0 : _GEN_1609; // @[CPU6502.scala 220:17 66:22]
  wire [7:0] _GEN_1629 = 8'hc8 == opcode ? regX : _GEN_1606; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_1630 = 8'hc8 == opcode ? regA : _GEN_1611; // @[CPU6502.scala 18:21 66:22]
  wire  _GEN_1631 = 8'hc8 == opcode ? flagC : _GEN_1612; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_1632 = 8'hc8 == opcode ? flagD : _GEN_1613; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_1633 = 8'hc8 == opcode ? flagI : _GEN_1614; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_1634 = 8'hc8 == opcode ? flagV : _GEN_1615; // @[CPU6502.scala 30:22 66:22]
  wire [15:0] _GEN_1635 = 8'hc8 == opcode ? regPC : _GEN_1616; // @[CPU6502.scala 42:14 66:22]
  wire  _GEN_1636 = 8'hc8 == opcode ? 1'h0 : _GEN_1617; // @[CPU6502.scala 45:14 66:22]
  wire [15:0] _GEN_1637 = 8'hc8 == opcode ? operand : _GEN_1618; // @[CPU6502.scala 66:22 38:24]
  wire [15:0] _GEN_1638 = 8'hc8 == opcode ? regPC : _GEN_1619; // @[CPU6502.scala 22:22 66:22]
  wire [2:0] _GEN_1639 = 8'hc8 == opcode ? cycle : _GEN_1620; // @[CPU6502.scala 39:22 66:22]
  wire [7:0] _GEN_1640 = 8'hc8 == opcode ? 8'h0 : _GEN_1621; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1641 = 8'hc8 == opcode ? 1'h0 : _GEN_1622; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_1642 = 8'hc8 == opcode ? regSP : _GEN_1623; // @[CPU6502.scala 21:22 66:22]
  wire [7:0] _GEN_1644 = 8'he8 == opcode ? result_3 : _GEN_1629; // @[CPU6502.scala 210:16 66:22]
  wire  _GEN_1645 = 8'he8 == opcode ? result_3[7] : _GEN_1626; // @[CPU6502.scala 50:11 66:22]
  wire  _GEN_1646 = 8'he8 == opcode ? result_3 == 8'h0 : _GEN_1627; // @[CPU6502.scala 51:11 66:22]
  wire [1:0] _GEN_1647 = 8'he8 == opcode ? 2'h0 : _GEN_1628; // @[CPU6502.scala 212:17 66:22]
  wire [7:0] _GEN_1648 = 8'he8 == opcode ? regY : _GEN_1625; // @[CPU6502.scala 20:21 66:22]
  wire [7:0] _GEN_1649 = 8'he8 == opcode ? regA : _GEN_1630; // @[CPU6502.scala 18:21 66:22]
  wire  _GEN_1650 = 8'he8 == opcode ? flagC : _GEN_1631; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_1651 = 8'he8 == opcode ? flagD : _GEN_1632; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_1652 = 8'he8 == opcode ? flagI : _GEN_1633; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_1653 = 8'he8 == opcode ? flagV : _GEN_1634; // @[CPU6502.scala 30:22 66:22]
  wire [15:0] _GEN_1654 = 8'he8 == opcode ? regPC : _GEN_1635; // @[CPU6502.scala 42:14 66:22]
  wire  _GEN_1655 = 8'he8 == opcode ? 1'h0 : _GEN_1636; // @[CPU6502.scala 45:14 66:22]
  wire [15:0] _GEN_1656 = 8'he8 == opcode ? operand : _GEN_1637; // @[CPU6502.scala 66:22 38:24]
  wire [15:0] _GEN_1657 = 8'he8 == opcode ? regPC : _GEN_1638; // @[CPU6502.scala 22:22 66:22]
  wire [2:0] _GEN_1658 = 8'he8 == opcode ? cycle : _GEN_1639; // @[CPU6502.scala 39:22 66:22]
  wire [7:0] _GEN_1659 = 8'he8 == opcode ? 8'h0 : _GEN_1640; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1660 = 8'he8 == opcode ? 1'h0 : _GEN_1641; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_1661 = 8'he8 == opcode ? regSP : _GEN_1642; // @[CPU6502.scala 21:22 66:22]
  wire [15:0] _GEN_1663 = 8'h49 == opcode ? regPC : _GEN_1654; // @[CPU6502.scala 66:22]
  wire  _GEN_1664 = 8'h49 == opcode ? _T_3 : _GEN_1655; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_1665 = 8'h49 == opcode ? _GEN_82 : _GEN_1649; // @[CPU6502.scala 66:22]
  wire  _GEN_1666 = 8'h49 == opcode ? _GEN_83 : _GEN_1645; // @[CPU6502.scala 66:22]
  wire  _GEN_1667 = 8'h49 == opcode ? _GEN_84 : _GEN_1646; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_1668 = 8'h49 == opcode ? _GEN_5 : _GEN_1657; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_1669 = 8'h49 == opcode ? _GEN_6 : _GEN_1647; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_1670 = 8'h49 == opcode ? regX : _GEN_1644; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_1671 = 8'h49 == opcode ? regY : _GEN_1648; // @[CPU6502.scala 20:21 66:22]
  wire  _GEN_1672 = 8'h49 == opcode ? flagC : _GEN_1650; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_1673 = 8'h49 == opcode ? flagD : _GEN_1651; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_1674 = 8'h49 == opcode ? flagI : _GEN_1652; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_1675 = 8'h49 == opcode ? flagV : _GEN_1653; // @[CPU6502.scala 30:22 66:22]
  wire [15:0] _GEN_1676 = 8'h49 == opcode ? operand : _GEN_1656; // @[CPU6502.scala 66:22 38:24]
  wire [2:0] _GEN_1677 = 8'h49 == opcode ? cycle : _GEN_1658; // @[CPU6502.scala 39:22 66:22]
  wire [7:0] _GEN_1678 = 8'h49 == opcode ? 8'h0 : _GEN_1659; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1679 = 8'h49 == opcode ? 1'h0 : _GEN_1660; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_1680 = 8'h49 == opcode ? regSP : _GEN_1661; // @[CPU6502.scala 21:22 66:22]
  wire [15:0] _GEN_1682 = 8'h9 == opcode ? regPC : _GEN_1663; // @[CPU6502.scala 66:22]
  wire  _GEN_1683 = 8'h9 == opcode ? _T_3 : _GEN_1664; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_1684 = 8'h9 == opcode ? _GEN_75 : _GEN_1665; // @[CPU6502.scala 66:22]
  wire  _GEN_1685 = 8'h9 == opcode ? _GEN_76 : _GEN_1666; // @[CPU6502.scala 66:22]
  wire  _GEN_1686 = 8'h9 == opcode ? _GEN_77 : _GEN_1667; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_1687 = 8'h9 == opcode ? _GEN_5 : _GEN_1668; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_1688 = 8'h9 == opcode ? _GEN_6 : _GEN_1669; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_1689 = 8'h9 == opcode ? regX : _GEN_1670; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_1690 = 8'h9 == opcode ? regY : _GEN_1671; // @[CPU6502.scala 20:21 66:22]
  wire  _GEN_1691 = 8'h9 == opcode ? flagC : _GEN_1672; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_1692 = 8'h9 == opcode ? flagD : _GEN_1673; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_1693 = 8'h9 == opcode ? flagI : _GEN_1674; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_1694 = 8'h9 == opcode ? flagV : _GEN_1675; // @[CPU6502.scala 30:22 66:22]
  wire [15:0] _GEN_1695 = 8'h9 == opcode ? operand : _GEN_1676; // @[CPU6502.scala 66:22 38:24]
  wire [2:0] _GEN_1696 = 8'h9 == opcode ? cycle : _GEN_1677; // @[CPU6502.scala 39:22 66:22]
  wire [7:0] _GEN_1697 = 8'h9 == opcode ? 8'h0 : _GEN_1678; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1698 = 8'h9 == opcode ? 1'h0 : _GEN_1679; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_1699 = 8'h9 == opcode ? regSP : _GEN_1680; // @[CPU6502.scala 21:22 66:22]
  wire [15:0] _GEN_1701 = 8'h29 == opcode ? regPC : _GEN_1682; // @[CPU6502.scala 66:22]
  wire  _GEN_1702 = 8'h29 == opcode ? _T_3 : _GEN_1683; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_1703 = 8'h29 == opcode ? _GEN_68 : _GEN_1684; // @[CPU6502.scala 66:22]
  wire  _GEN_1704 = 8'h29 == opcode ? _GEN_69 : _GEN_1685; // @[CPU6502.scala 66:22]
  wire  _GEN_1705 = 8'h29 == opcode ? _GEN_70 : _GEN_1686; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_1706 = 8'h29 == opcode ? _GEN_5 : _GEN_1687; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_1707 = 8'h29 == opcode ? _GEN_6 : _GEN_1688; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_1708 = 8'h29 == opcode ? regX : _GEN_1689; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_1709 = 8'h29 == opcode ? regY : _GEN_1690; // @[CPU6502.scala 20:21 66:22]
  wire  _GEN_1710 = 8'h29 == opcode ? flagC : _GEN_1691; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_1711 = 8'h29 == opcode ? flagD : _GEN_1692; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_1712 = 8'h29 == opcode ? flagI : _GEN_1693; // @[CPU6502.scala 27:22 66:22]
  wire  _GEN_1713 = 8'h29 == opcode ? flagV : _GEN_1694; // @[CPU6502.scala 30:22 66:22]
  wire [15:0] _GEN_1714 = 8'h29 == opcode ? operand : _GEN_1695; // @[CPU6502.scala 66:22 38:24]
  wire [2:0] _GEN_1715 = 8'h29 == opcode ? cycle : _GEN_1696; // @[CPU6502.scala 39:22 66:22]
  wire [7:0] _GEN_1716 = 8'h29 == opcode ? 8'h0 : _GEN_1697; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1717 = 8'h29 == opcode ? 1'h0 : _GEN_1698; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_1718 = 8'h29 == opcode ? regSP : _GEN_1699; // @[CPU6502.scala 21:22 66:22]
  wire [15:0] _GEN_1720 = 8'he9 == opcode ? regPC : _GEN_1701; // @[CPU6502.scala 66:22]
  wire  _GEN_1721 = 8'he9 == opcode ? _T_3 : _GEN_1702; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_1722 = 8'he9 == opcode ? _GEN_59 : _GEN_1703; // @[CPU6502.scala 66:22]
  wire  _GEN_1723 = 8'he9 == opcode ? _GEN_60 : _GEN_1710; // @[CPU6502.scala 66:22]
  wire  _GEN_1724 = 8'he9 == opcode ? _GEN_61 : _GEN_1704; // @[CPU6502.scala 66:22]
  wire  _GEN_1725 = 8'he9 == opcode ? _GEN_62 : _GEN_1705; // @[CPU6502.scala 66:22]
  wire  _GEN_1726 = 8'he9 == opcode ? _GEN_63 : _GEN_1713; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_1727 = 8'he9 == opcode ? _GEN_5 : _GEN_1706; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_1728 = 8'he9 == opcode ? _GEN_6 : _GEN_1707; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_1729 = 8'he9 == opcode ? regX : _GEN_1708; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_1730 = 8'he9 == opcode ? regY : _GEN_1709; // @[CPU6502.scala 20:21 66:22]
  wire  _GEN_1731 = 8'he9 == opcode ? flagD : _GEN_1711; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_1732 = 8'he9 == opcode ? flagI : _GEN_1712; // @[CPU6502.scala 27:22 66:22]
  wire [15:0] _GEN_1733 = 8'he9 == opcode ? operand : _GEN_1714; // @[CPU6502.scala 66:22 38:24]
  wire [2:0] _GEN_1734 = 8'he9 == opcode ? cycle : _GEN_1715; // @[CPU6502.scala 39:22 66:22]
  wire [7:0] _GEN_1735 = 8'he9 == opcode ? 8'h0 : _GEN_1716; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1736 = 8'he9 == opcode ? 1'h0 : _GEN_1717; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_1737 = 8'he9 == opcode ? regSP : _GEN_1718; // @[CPU6502.scala 21:22 66:22]
  wire [15:0] _GEN_1739 = 8'h69 == opcode ? regPC : _GEN_1720; // @[CPU6502.scala 66:22]
  wire  _GEN_1740 = 8'h69 == opcode ? _T_3 : _GEN_1721; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_1741 = 8'h69 == opcode ? _GEN_50 : _GEN_1722; // @[CPU6502.scala 66:22]
  wire  _GEN_1742 = 8'h69 == opcode ? _GEN_51 : _GEN_1723; // @[CPU6502.scala 66:22]
  wire  _GEN_1743 = 8'h69 == opcode ? _GEN_52 : _GEN_1724; // @[CPU6502.scala 66:22]
  wire  _GEN_1744 = 8'h69 == opcode ? _GEN_53 : _GEN_1725; // @[CPU6502.scala 66:22]
  wire  _GEN_1745 = 8'h69 == opcode ? _GEN_54 : _GEN_1726; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_1746 = 8'h69 == opcode ? _GEN_5 : _GEN_1727; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_1747 = 8'h69 == opcode ? _GEN_6 : _GEN_1728; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_1748 = 8'h69 == opcode ? regX : _GEN_1729; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_1749 = 8'h69 == opcode ? regY : _GEN_1730; // @[CPU6502.scala 20:21 66:22]
  wire  _GEN_1750 = 8'h69 == opcode ? flagD : _GEN_1731; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_1751 = 8'h69 == opcode ? flagI : _GEN_1732; // @[CPU6502.scala 27:22 66:22]
  wire [15:0] _GEN_1752 = 8'h69 == opcode ? operand : _GEN_1733; // @[CPU6502.scala 66:22 38:24]
  wire [2:0] _GEN_1753 = 8'h69 == opcode ? cycle : _GEN_1734; // @[CPU6502.scala 39:22 66:22]
  wire [7:0] _GEN_1754 = 8'h69 == opcode ? 8'h0 : _GEN_1735; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1755 = 8'h69 == opcode ? 1'h0 : _GEN_1736; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_1756 = 8'h69 == opcode ? regSP : _GEN_1737; // @[CPU6502.scala 21:22 66:22]
  wire [15:0] _GEN_1758 = 8'h85 == opcode ? _GEN_13 : _GEN_1739; // @[CPU6502.scala 66:22]
  wire  _GEN_1759 = 8'h85 == opcode ? _T_3 : _GEN_1740; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_1760 = 8'h85 == opcode ? _GEN_15 : _GEN_1752; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_1761 = 8'h85 == opcode ? _GEN_5 : _GEN_1746; // @[CPU6502.scala 66:22]
  wire [2:0] _GEN_1762 = 8'h85 == opcode ? _GEN_17 : _GEN_1753; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_1763 = 8'h85 == opcode ? _GEN_45 : _GEN_1754; // @[CPU6502.scala 66:22]
  wire  _GEN_1764 = 8'h85 == opcode ? _GEN_46 : _GEN_1755; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_1765 = 8'h85 == opcode ? _GEN_21 : _GEN_1747; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_1766 = 8'h85 == opcode ? regA : _GEN_1741; // @[CPU6502.scala 18:21 66:22]
  wire  _GEN_1767 = 8'h85 == opcode ? flagC : _GEN_1742; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_1768 = 8'h85 == opcode ? flagN : _GEN_1743; // @[CPU6502.scala 31:22 66:22]
  wire  _GEN_1769 = 8'h85 == opcode ? flagZ : _GEN_1744; // @[CPU6502.scala 26:22 66:22]
  wire  _GEN_1770 = 8'h85 == opcode ? flagV : _GEN_1745; // @[CPU6502.scala 30:22 66:22]
  wire [7:0] _GEN_1771 = 8'h85 == opcode ? regX : _GEN_1748; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_1772 = 8'h85 == opcode ? regY : _GEN_1749; // @[CPU6502.scala 20:21 66:22]
  wire  _GEN_1773 = 8'h85 == opcode ? flagD : _GEN_1750; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_1774 = 8'h85 == opcode ? flagI : _GEN_1751; // @[CPU6502.scala 27:22 66:22]
  wire [7:0] _GEN_1775 = 8'h85 == opcode ? regSP : _GEN_1756; // @[CPU6502.scala 21:22 66:22]
  wire [15:0] _GEN_1777 = 8'ha0 == opcode ? regPC : _GEN_1758; // @[CPU6502.scala 66:22]
  wire  _GEN_1778 = 8'ha0 == opcode ? _T_3 : _GEN_1759; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_1779 = 8'ha0 == opcode ? _GEN_31 : _GEN_1772; // @[CPU6502.scala 66:22]
  wire  _GEN_1780 = 8'ha0 == opcode ? _GEN_3 : _GEN_1768; // @[CPU6502.scala 66:22]
  wire  _GEN_1781 = 8'ha0 == opcode ? _GEN_4 : _GEN_1769; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_1782 = 8'ha0 == opcode ? _GEN_5 : _GEN_1761; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_1783 = 8'ha0 == opcode ? _GEN_6 : _GEN_1765; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_1784 = 8'ha0 == opcode ? operand : _GEN_1760; // @[CPU6502.scala 66:22 38:24]
  wire [2:0] _GEN_1785 = 8'ha0 == opcode ? cycle : _GEN_1762; // @[CPU6502.scala 39:22 66:22]
  wire [7:0] _GEN_1786 = 8'ha0 == opcode ? 8'h0 : _GEN_1763; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1787 = 8'ha0 == opcode ? 1'h0 : _GEN_1764; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_1788 = 8'ha0 == opcode ? regA : _GEN_1766; // @[CPU6502.scala 18:21 66:22]
  wire  _GEN_1789 = 8'ha0 == opcode ? flagC : _GEN_1767; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_1790 = 8'ha0 == opcode ? flagV : _GEN_1770; // @[CPU6502.scala 30:22 66:22]
  wire [7:0] _GEN_1791 = 8'ha0 == opcode ? regX : _GEN_1771; // @[CPU6502.scala 19:21 66:22]
  wire  _GEN_1792 = 8'ha0 == opcode ? flagD : _GEN_1773; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_1793 = 8'ha0 == opcode ? flagI : _GEN_1774; // @[CPU6502.scala 27:22 66:22]
  wire [7:0] _GEN_1794 = 8'ha0 == opcode ? regSP : _GEN_1775; // @[CPU6502.scala 21:22 66:22]
  wire [15:0] _GEN_1796 = 8'ha2 == opcode ? regPC : _GEN_1777; // @[CPU6502.scala 66:22]
  wire  _GEN_1797 = 8'ha2 == opcode ? _T_3 : _GEN_1778; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_1798 = 8'ha2 == opcode ? _GEN_24 : _GEN_1791; // @[CPU6502.scala 66:22]
  wire  _GEN_1799 = 8'ha2 == opcode ? _GEN_3 : _GEN_1780; // @[CPU6502.scala 66:22]
  wire  _GEN_1800 = 8'ha2 == opcode ? _GEN_4 : _GEN_1781; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_1801 = 8'ha2 == opcode ? _GEN_5 : _GEN_1782; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_1802 = 8'ha2 == opcode ? _GEN_6 : _GEN_1783; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_1803 = 8'ha2 == opcode ? regY : _GEN_1779; // @[CPU6502.scala 20:21 66:22]
  wire [15:0] _GEN_1804 = 8'ha2 == opcode ? operand : _GEN_1784; // @[CPU6502.scala 66:22 38:24]
  wire [2:0] _GEN_1805 = 8'ha2 == opcode ? cycle : _GEN_1785; // @[CPU6502.scala 39:22 66:22]
  wire [7:0] _GEN_1806 = 8'ha2 == opcode ? 8'h0 : _GEN_1786; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1807 = 8'ha2 == opcode ? 1'h0 : _GEN_1787; // @[CPU6502.scala 44:15 66:22]
  wire [7:0] _GEN_1808 = 8'ha2 == opcode ? regA : _GEN_1788; // @[CPU6502.scala 18:21 66:22]
  wire  _GEN_1809 = 8'ha2 == opcode ? flagC : _GEN_1789; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_1810 = 8'ha2 == opcode ? flagV : _GEN_1790; // @[CPU6502.scala 30:22 66:22]
  wire  _GEN_1811 = 8'ha2 == opcode ? flagD : _GEN_1792; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_1812 = 8'ha2 == opcode ? flagI : _GEN_1793; // @[CPU6502.scala 27:22 66:22]
  wire [7:0] _GEN_1813 = 8'ha2 == opcode ? regSP : _GEN_1794; // @[CPU6502.scala 21:22 66:22]
  wire [15:0] _GEN_1815 = 8'ha5 == opcode ? _GEN_13 : _GEN_1796; // @[CPU6502.scala 66:22]
  wire  _GEN_1816 = 8'ha5 == opcode ? _GEN_14 : _GEN_1797; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_1817 = 8'ha5 == opcode ? _GEN_15 : _GEN_1804; // @[CPU6502.scala 66:22]
  wire [15:0] _GEN_1818 = 8'ha5 == opcode ? _GEN_5 : _GEN_1801; // @[CPU6502.scala 66:22]
  wire [2:0] _GEN_1819 = 8'ha5 == opcode ? _GEN_17 : _GEN_1805; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_1820 = 8'ha5 == opcode ? _GEN_18 : _GEN_1808; // @[CPU6502.scala 66:22]
  wire  _GEN_1821 = 8'ha5 == opcode ? _GEN_19 : _GEN_1799; // @[CPU6502.scala 66:22]
  wire  _GEN_1822 = 8'ha5 == opcode ? _GEN_20 : _GEN_1800; // @[CPU6502.scala 66:22]
  wire [1:0] _GEN_1823 = 8'ha5 == opcode ? _GEN_21 : _GEN_1802; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_1824 = 8'ha5 == opcode ? regX : _GEN_1798; // @[CPU6502.scala 19:21 66:22]
  wire [7:0] _GEN_1825 = 8'ha5 == opcode ? regY : _GEN_1803; // @[CPU6502.scala 20:21 66:22]
  wire [7:0] _GEN_1826 = 8'ha5 == opcode ? 8'h0 : _GEN_1806; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1827 = 8'ha5 == opcode ? 1'h0 : _GEN_1807; // @[CPU6502.scala 44:15 66:22]
  wire  _GEN_1828 = 8'ha5 == opcode ? flagC : _GEN_1809; // @[CPU6502.scala 25:22 66:22]
  wire  _GEN_1829 = 8'ha5 == opcode ? flagV : _GEN_1810; // @[CPU6502.scala 30:22 66:22]
  wire  _GEN_1830 = 8'ha5 == opcode ? flagD : _GEN_1811; // @[CPU6502.scala 28:22 66:22]
  wire  _GEN_1831 = 8'ha5 == opcode ? flagI : _GEN_1812; // @[CPU6502.scala 27:22 66:22]
  wire [7:0] _GEN_1832 = 8'ha5 == opcode ? regSP : _GEN_1813; // @[CPU6502.scala 21:22 66:22]
  wire [15:0] _GEN_1834 = 8'ha9 == opcode ? regPC : _GEN_1815; // @[CPU6502.scala 66:22]
  wire  _GEN_1835 = 8'ha9 == opcode ? _T_3 : _GEN_1816; // @[CPU6502.scala 66:22]
  wire [7:0] _GEN_1845 = 8'ha9 == opcode ? 8'h0 : _GEN_1826; // @[CPU6502.scala 43:17 66:22]
  wire  _GEN_1846 = 8'ha9 == opcode ? 1'h0 : _GEN_1827; // @[CPU6502.scala 44:15 66:22]
  wire [15:0] _GEN_1853 = 2'h1 == state ? _GEN_1834 : regPC; // @[CPU6502.scala 42:14 55:17]
  wire  _GEN_1854 = 2'h1 == state & _GEN_1835; // @[CPU6502.scala 45:14 55:17]
  wire [7:0] _GEN_1864 = 2'h1 == state ? _GEN_1845 : 8'h0; // @[CPU6502.scala 43:17 55:17]
  assign io_memAddr = 2'h0 == state ? regPC : _GEN_1853; // @[CPU6502.scala 55:17 57:18]
  assign io_memDataOut = 2'h0 == state ? 8'h0 : _GEN_1864; // @[CPU6502.scala 43:17 55:17]
  assign io_memWrite = 2'h0 == state ? 1'h0 : 2'h1 == state & _GEN_1846; // @[CPU6502.scala 44:15 55:17]
  assign io_memRead = 2'h0 == state | _GEN_1854; // @[CPU6502.scala 55:17 58:18]
  assign io_debug_regA = regA; // @[CPU6502.scala 1076:17]
  assign io_debug_regX = regX; // @[CPU6502.scala 1077:17]
  assign io_debug_regY = regY; // @[CPU6502.scala 1078:17]
  assign io_debug_regPC = regPC; // @[CPU6502.scala 1079:18]
  assign io_debug_regSP = regSP; // @[CPU6502.scala 1080:18]
  assign io_debug_flagC = flagC; // @[CPU6502.scala 1081:18]
  assign io_debug_flagZ = flagZ; // @[CPU6502.scala 1082:18]
  assign io_debug_flagN = flagN; // @[CPU6502.scala 1083:18]
  assign io_debug_flagV = flagV; // @[CPU6502.scala 1084:18]
  assign io_debug_opcode = opcode; // @[CPU6502.scala 1085:19]
  always @(posedge clock) begin
    if (reset) begin // @[CPU6502.scala 18:21]
      regA <= 8'h0; // @[CPU6502.scala 18:21]
    end else if (!(2'h0 == state)) begin // @[CPU6502.scala 55:17]
      if (2'h1 == state) begin // @[CPU6502.scala 55:17]
        if (8'ha9 == opcode) begin // @[CPU6502.scala 66:22]
          regA <= _GEN_2;
        end else begin
          regA <= _GEN_1820;
        end
      end
    end
    if (reset) begin // @[CPU6502.scala 19:21]
      regX <= 8'h0; // @[CPU6502.scala 19:21]
    end else if (!(2'h0 == state)) begin // @[CPU6502.scala 55:17]
      if (2'h1 == state) begin // @[CPU6502.scala 55:17]
        if (!(8'ha9 == opcode)) begin // @[CPU6502.scala 66:22]
          regX <= _GEN_1824;
        end
      end
    end
    if (reset) begin // @[CPU6502.scala 20:21]
      regY <= 8'h0; // @[CPU6502.scala 20:21]
    end else if (!(2'h0 == state)) begin // @[CPU6502.scala 55:17]
      if (2'h1 == state) begin // @[CPU6502.scala 55:17]
        if (!(8'ha9 == opcode)) begin // @[CPU6502.scala 66:22]
          regY <= _GEN_1825;
        end
      end
    end
    if (reset) begin // @[CPU6502.scala 21:22]
      regSP <= 8'hff; // @[CPU6502.scala 21:22]
    end else if (!(2'h0 == state)) begin // @[CPU6502.scala 55:17]
      if (2'h1 == state) begin // @[CPU6502.scala 55:17]
        if (!(8'ha9 == opcode)) begin // @[CPU6502.scala 66:22]
          regSP <= _GEN_1832;
        end
      end
    end
    if (reset) begin // @[CPU6502.scala 22:22]
      regPC <= 16'h0; // @[CPU6502.scala 22:22]
    end else if (2'h0 == state) begin // @[CPU6502.scala 55:17]
      regPC <= _regPC_T_1; // @[CPU6502.scala 60:13]
    end else if (2'h1 == state) begin // @[CPU6502.scala 55:17]
      if (8'ha9 == opcode) begin // @[CPU6502.scala 66:22]
        regPC <= _GEN_5;
      end else begin
        regPC <= _GEN_1818;
      end
    end
    if (reset) begin // @[CPU6502.scala 25:22]
      flagC <= 1'h0; // @[CPU6502.scala 25:22]
    end else if (!(2'h0 == state)) begin // @[CPU6502.scala 55:17]
      if (2'h1 == state) begin // @[CPU6502.scala 55:17]
        if (!(8'ha9 == opcode)) begin // @[CPU6502.scala 66:22]
          flagC <= _GEN_1828;
        end
      end
    end
    if (reset) begin // @[CPU6502.scala 26:22]
      flagZ <= 1'h0; // @[CPU6502.scala 26:22]
    end else if (!(2'h0 == state)) begin // @[CPU6502.scala 55:17]
      if (2'h1 == state) begin // @[CPU6502.scala 55:17]
        if (8'ha9 == opcode) begin // @[CPU6502.scala 66:22]
          flagZ <= _GEN_4;
        end else begin
          flagZ <= _GEN_1822;
        end
      end
    end
    if (reset) begin // @[CPU6502.scala 27:22]
      flagI <= 1'h0; // @[CPU6502.scala 27:22]
    end else if (!(2'h0 == state)) begin // @[CPU6502.scala 55:17]
      if (2'h1 == state) begin // @[CPU6502.scala 55:17]
        if (!(8'ha9 == opcode)) begin // @[CPU6502.scala 66:22]
          flagI <= _GEN_1831;
        end
      end
    end
    if (reset) begin // @[CPU6502.scala 28:22]
      flagD <= 1'h0; // @[CPU6502.scala 28:22]
    end else if (!(2'h0 == state)) begin // @[CPU6502.scala 55:17]
      if (2'h1 == state) begin // @[CPU6502.scala 55:17]
        if (!(8'ha9 == opcode)) begin // @[CPU6502.scala 66:22]
          flagD <= _GEN_1830;
        end
      end
    end
    if (reset) begin // @[CPU6502.scala 30:22]
      flagV <= 1'h0; // @[CPU6502.scala 30:22]
    end else if (!(2'h0 == state)) begin // @[CPU6502.scala 55:17]
      if (2'h1 == state) begin // @[CPU6502.scala 55:17]
        if (!(8'ha9 == opcode)) begin // @[CPU6502.scala 66:22]
          flagV <= _GEN_1829;
        end
      end
    end
    if (reset) begin // @[CPU6502.scala 31:22]
      flagN <= 1'h0; // @[CPU6502.scala 31:22]
    end else if (!(2'h0 == state)) begin // @[CPU6502.scala 55:17]
      if (2'h1 == state) begin // @[CPU6502.scala 55:17]
        if (8'ha9 == opcode) begin // @[CPU6502.scala 66:22]
          flagN <= _GEN_3;
        end else begin
          flagN <= _GEN_1821;
        end
      end
    end
    if (reset) begin // @[CPU6502.scala 35:22]
      state <= 2'h0; // @[CPU6502.scala 35:22]
    end else if (2'h0 == state) begin // @[CPU6502.scala 55:17]
      state <= 2'h1; // @[CPU6502.scala 61:13]
    end else if (2'h1 == state) begin // @[CPU6502.scala 55:17]
      if (8'ha9 == opcode) begin // @[CPU6502.scala 66:22]
        state <= _GEN_6;
      end else begin
        state <= _GEN_1823;
      end
    end
    if (reset) begin // @[CPU6502.scala 37:23]
      opcode <= 8'h0; // @[CPU6502.scala 37:23]
    end else if (2'h0 == state) begin // @[CPU6502.scala 55:17]
      opcode <= io_memDataIn; // @[CPU6502.scala 59:14]
    end
    if (reset) begin // @[CPU6502.scala 38:24]
      operand <= 16'h0; // @[CPU6502.scala 38:24]
    end else if (!(2'h0 == state)) begin // @[CPU6502.scala 55:17]
      if (2'h1 == state) begin // @[CPU6502.scala 55:17]
        if (!(8'ha9 == opcode)) begin // @[CPU6502.scala 66:22]
          operand <= _GEN_1817;
        end
      end
    end
    if (reset) begin // @[CPU6502.scala 39:22]
      cycle <= 3'h0; // @[CPU6502.scala 39:22]
    end else if (!(2'h0 == state)) begin // @[CPU6502.scala 55:17]
      if (2'h1 == state) begin // @[CPU6502.scala 55:17]
        if (!(8'ha9 == opcode)) begin // @[CPU6502.scala 66:22]
          cycle <= _GEN_1819;
        end
      end
    end
  end
endmodule
module PPU(
  input        clock,
  input        reset,
  input  [2:0] io_cpuAddr,
  input  [7:0] io_cpuDataIn,
  output [7:0] io_cpuDataOut,
  input        io_cpuWrite,
  input        io_cpuRead,
  output [8:0] io_pixelX,
  output [8:0] io_pixelY,
  output       io_vblank
);
  reg [7:0] vram [0:2047]; // @[PPU.scala 47:25]
  wire  vram_io_cpuDataOut_MPORT_1_en; // @[PPU.scala 47:25]
  wire [10:0] vram_io_cpuDataOut_MPORT_1_addr; // @[PPU.scala 47:25]
  wire [7:0] vram_io_cpuDataOut_MPORT_1_data; // @[PPU.scala 47:25]
  wire [7:0] vram_MPORT_1_data; // @[PPU.scala 47:25]
  wire [10:0] vram_MPORT_1_addr; // @[PPU.scala 47:25]
  wire  vram_MPORT_1_mask; // @[PPU.scala 47:25]
  wire  vram_MPORT_1_en; // @[PPU.scala 47:25]
  reg  vram_io_cpuDataOut_MPORT_1_en_pipe_0;
  reg [10:0] vram_io_cpuDataOut_MPORT_1_addr_pipe_0;
  reg [7:0] oam [0:255]; // @[PPU.scala 48:24]
  wire  oam_io_cpuDataOut_MPORT_en; // @[PPU.scala 48:24]
  wire [7:0] oam_io_cpuDataOut_MPORT_addr; // @[PPU.scala 48:24]
  wire [7:0] oam_io_cpuDataOut_MPORT_data; // @[PPU.scala 48:24]
  wire [7:0] oam_MPORT_data; // @[PPU.scala 48:24]
  wire [7:0] oam_MPORT_addr; // @[PPU.scala 48:24]
  wire  oam_MPORT_mask; // @[PPU.scala 48:24]
  wire  oam_MPORT_en; // @[PPU.scala 48:24]
  reg  oam_io_cpuDataOut_MPORT_en_pipe_0;
  reg [7:0] oam_io_cpuDataOut_MPORT_addr_pipe_0;
  reg [7:0] oamAddr; // @[PPU.scala 40:24]
  reg  ppuAddrLatch; // @[PPU.scala 43:29]
  reg [15:0] ppuAddrReg; // @[PPU.scala 44:27]
  reg [8:0] scanlineX; // @[PPU.scala 52:26]
  reg [8:0] scanlineY; // @[PPU.scala 53:26]
  reg  vblankFlag; // @[PPU.scala 56:27]
  wire [8:0] _scanlineX_T_1 = scanlineX + 9'h1; // @[PPU.scala 60:26]
  wire [8:0] _scanlineY_T_1 = scanlineY + 9'h1; // @[PPU.scala 63:28]
  wire  _T_1 = scanlineY == 9'h105; // @[PPU.scala 65:20]
  wire  _T_3 = scanlineX == 9'h1; // @[PPU.scala 71:41]
  wire  _GEN_4 = scanlineY == 9'hf1 & scanlineX == 9'h1 | vblankFlag; // @[PPU.scala 71:50 72:16 56:27]
  wire  _GEN_6 = _T_1 & _T_3 ? 1'h0 : _GEN_4; // @[PPU.scala 78:50 79:16]
  wire [7:0] _io_cpuDataOut_T = {vblankFlag,7'h0}; // @[Cat.scala 33:92]
  wire  _T_10 = 3'h4 == io_cpuAddr; // @[PPU.scala 87:24]
  wire  _T_11 = 3'h7 == io_cpuAddr; // @[PPU.scala 87:24]
  wire [15:0] _ppuAddrReg_T_1 = ppuAddrReg + 16'h1; // @[PPU.scala 99:34]
  wire [7:0] _GEN_17 = 3'h7 == io_cpuAddr ? vram_io_cpuDataOut_MPORT_1_data : 8'h0; // @[PPU.scala 84:17 87:24 98:23]
  wire [15:0] _GEN_18 = 3'h7 == io_cpuAddr ? _ppuAddrReg_T_1 : ppuAddrReg; // @[PPU.scala 87:24 99:20 44:27]
  wire [7:0] _GEN_22 = 3'h4 == io_cpuAddr ? oam_io_cpuDataOut_MPORT_data : _GEN_17; // @[PPU.scala 87:24 94:23]
  wire  _GEN_23 = 3'h4 == io_cpuAddr ? 1'h0 : 3'h7 == io_cpuAddr; // @[PPU.scala 87:24 47:25]
  wire [15:0] _GEN_26 = 3'h4 == io_cpuAddr ? ppuAddrReg : _GEN_18; // @[PPU.scala 87:24 44:27]
  wire [7:0] _GEN_27 = 3'h2 == io_cpuAddr ? _io_cpuDataOut_T : _GEN_22; // @[PPU.scala 87:24 89:23]
  wire  _GEN_29 = 3'h2 == io_cpuAddr ? 1'h0 : ppuAddrLatch; // @[PPU.scala 87:24 91:22 43:29]
  wire  _GEN_30 = 3'h2 == io_cpuAddr ? 1'h0 : 3'h4 == io_cpuAddr; // @[PPU.scala 48:24 87:24]
  wire  _GEN_33 = 3'h2 == io_cpuAddr ? 1'h0 : _GEN_23; // @[PPU.scala 87:24 47:25]
  wire [15:0] _GEN_36 = 3'h2 == io_cpuAddr ? ppuAddrReg : _GEN_26; // @[PPU.scala 87:24 44:27]
  wire  _GEN_39 = io_cpuRead ? _GEN_29 : ppuAddrLatch; // @[PPU.scala 86:20 43:29]
  wire [15:0] _GEN_46 = io_cpuRead ? _GEN_36 : ppuAddrReg; // @[PPU.scala 86:20 44:27]
  wire [7:0] _oamAddr_T_1 = oamAddr + 8'h1; // @[PPU.scala 117:28]
  wire  _T_17 = ~ppuAddrLatch; // @[PPU.scala 120:14]
  wire [13:0] _ppuAddrReg_T_3 = {io_cpuDataIn[5:0],8'h0}; // @[Cat.scala 33:92]
  wire [15:0] _ppuAddrReg_T_5 = {ppuAddrReg[15:8],io_cpuDataIn}; // @[Cat.scala 33:92]
  wire [15:0] _GEN_49 = _T_17 ? {{2'd0}, _ppuAddrReg_T_3} : _ppuAddrReg_T_5; // @[PPU.scala 128:29 129:22 131:22]
  wire [15:0] _GEN_55 = _T_11 ? _ppuAddrReg_T_1 : _GEN_46; // @[PPU.scala 105:24 138:20]
  wire [15:0] _GEN_56 = 3'h6 == io_cpuAddr ? _GEN_49 : _GEN_55; // @[PPU.scala 105:24]
  wire  _GEN_57 = 3'h6 == io_cpuAddr ? _T_17 : _GEN_39; // @[PPU.scala 105:24 133:22]
  wire  _GEN_60 = 3'h6 == io_cpuAddr ? 1'h0 : _T_11; // @[PPU.scala 105:24 47:25]
  wire  _GEN_65 = 3'h5 == io_cpuAddr ? _T_17 : _GEN_57; // @[PPU.scala 105:24 125:22]
  wire [15:0] _GEN_66 = 3'h5 == io_cpuAddr ? _GEN_46 : _GEN_56; // @[PPU.scala 105:24]
  wire  _GEN_69 = 3'h5 == io_cpuAddr ? 1'h0 : _GEN_60; // @[PPU.scala 105:24 47:25]
  wire [7:0] _GEN_77 = _T_10 ? _oamAddr_T_1 : oamAddr; // @[PPU.scala 105:24 117:17 40:24]
  wire  _GEN_80 = _T_10 ? _GEN_39 : _GEN_65; // @[PPU.scala 105:24]
  wire [15:0] _GEN_81 = _T_10 ? _GEN_46 : _GEN_66; // @[PPU.scala 105:24]
  wire  _GEN_84 = _T_10 ? 1'h0 : _GEN_69; // @[PPU.scala 105:24 47:25]
  wire [7:0] _GEN_87 = 3'h3 == io_cpuAddr ? io_cpuDataIn : _GEN_77; // @[PPU.scala 105:24 113:17]
  wire  _GEN_90 = 3'h3 == io_cpuAddr ? 1'h0 : _T_10; // @[PPU.scala 105:24 48:24]
  wire  _GEN_95 = 3'h3 == io_cpuAddr ? _GEN_39 : _GEN_80; // @[PPU.scala 105:24]
  wire [15:0] _GEN_96 = 3'h3 == io_cpuAddr ? _GEN_46 : _GEN_81; // @[PPU.scala 105:24]
  wire  _GEN_99 = 3'h3 == io_cpuAddr ? 1'h0 : _GEN_84; // @[PPU.scala 105:24 47:25]
  wire  _GEN_106 = 3'h1 == io_cpuAddr ? 1'h0 : _GEN_90; // @[PPU.scala 105:24 48:24]
  wire  _GEN_115 = 3'h1 == io_cpuAddr ? 1'h0 : _GEN_99; // @[PPU.scala 105:24 47:25]
  wire  _GEN_123 = 3'h0 == io_cpuAddr ? 1'h0 : _GEN_106; // @[PPU.scala 105:24 48:24]
  wire  _GEN_132 = 3'h0 == io_cpuAddr ? 1'h0 : _GEN_115; // @[PPU.scala 105:24 47:25]
  assign vram_io_cpuDataOut_MPORT_1_en = vram_io_cpuDataOut_MPORT_1_en_pipe_0;
  assign vram_io_cpuDataOut_MPORT_1_addr = vram_io_cpuDataOut_MPORT_1_addr_pipe_0;
  assign vram_io_cpuDataOut_MPORT_1_data = vram[vram_io_cpuDataOut_MPORT_1_addr]; // @[PPU.scala 47:25]
  assign vram_MPORT_1_data = io_cpuDataIn;
  assign vram_MPORT_1_addr = ppuAddrReg[10:0];
  assign vram_MPORT_1_mask = 1'h1;
  assign vram_MPORT_1_en = io_cpuWrite & _GEN_132;
  assign oam_io_cpuDataOut_MPORT_en = oam_io_cpuDataOut_MPORT_en_pipe_0;
  assign oam_io_cpuDataOut_MPORT_addr = oam_io_cpuDataOut_MPORT_addr_pipe_0;
  assign oam_io_cpuDataOut_MPORT_data = oam[oam_io_cpuDataOut_MPORT_addr]; // @[PPU.scala 48:24]
  assign oam_MPORT_data = io_cpuDataIn;
  assign oam_MPORT_addr = oamAddr;
  assign oam_MPORT_mask = 1'h1;
  assign oam_MPORT_en = io_cpuWrite & _GEN_123;
  assign io_cpuDataOut = io_cpuRead ? _GEN_27 : 8'h0; // @[PPU.scala 84:17 86:20]
  assign io_pixelX = scanlineX; // @[PPU.scala 144:13]
  assign io_pixelY = scanlineY; // @[PPU.scala 145:13]
  assign io_vblank = vblankFlag; // @[PPU.scala 147:13]
  always @(posedge clock) begin
    if (vram_MPORT_1_en & vram_MPORT_1_mask) begin
      vram[vram_MPORT_1_addr] <= vram_MPORT_1_data; // @[PPU.scala 47:25]
    end
    vram_io_cpuDataOut_MPORT_1_en_pipe_0 <= io_cpuRead & _GEN_33;
    if (io_cpuRead & _GEN_33) begin
      vram_io_cpuDataOut_MPORT_1_addr_pipe_0 <= ppuAddrReg[10:0];
    end
    if (oam_MPORT_en & oam_MPORT_mask) begin
      oam[oam_MPORT_addr] <= oam_MPORT_data; // @[PPU.scala 48:24]
    end
    oam_io_cpuDataOut_MPORT_en_pipe_0 <= io_cpuRead & _GEN_30;
    if (io_cpuRead & _GEN_30) begin
      oam_io_cpuDataOut_MPORT_addr_pipe_0 <= oamAddr;
    end
    if (reset) begin // @[PPU.scala 40:24]
      oamAddr <= 8'h0; // @[PPU.scala 40:24]
    end else if (io_cpuWrite) begin // @[PPU.scala 104:21]
      if (!(3'h0 == io_cpuAddr)) begin // @[PPU.scala 105:24]
        if (!(3'h1 == io_cpuAddr)) begin // @[PPU.scala 105:24]
          oamAddr <= _GEN_87;
        end
      end
    end
    if (reset) begin // @[PPU.scala 43:29]
      ppuAddrLatch <= 1'h0; // @[PPU.scala 43:29]
    end else if (io_cpuWrite) begin // @[PPU.scala 104:21]
      if (3'h0 == io_cpuAddr) begin // @[PPU.scala 105:24]
        ppuAddrLatch <= _GEN_39;
      end else if (3'h1 == io_cpuAddr) begin // @[PPU.scala 105:24]
        ppuAddrLatch <= _GEN_39;
      end else begin
        ppuAddrLatch <= _GEN_95;
      end
    end else begin
      ppuAddrLatch <= _GEN_39;
    end
    if (reset) begin // @[PPU.scala 44:27]
      ppuAddrReg <= 16'h0; // @[PPU.scala 44:27]
    end else if (io_cpuWrite) begin // @[PPU.scala 104:21]
      if (3'h0 == io_cpuAddr) begin // @[PPU.scala 105:24]
        ppuAddrReg <= _GEN_46;
      end else if (3'h1 == io_cpuAddr) begin // @[PPU.scala 105:24]
        ppuAddrReg <= _GEN_46;
      end else begin
        ppuAddrReg <= _GEN_96;
      end
    end else begin
      ppuAddrReg <= _GEN_46;
    end
    if (reset) begin // @[PPU.scala 52:26]
      scanlineX <= 9'h0; // @[PPU.scala 52:26]
    end else if (scanlineX == 9'h154) begin // @[PPU.scala 61:29]
      scanlineX <= 9'h0; // @[PPU.scala 62:15]
    end else begin
      scanlineX <= _scanlineX_T_1; // @[PPU.scala 60:13]
    end
    if (reset) begin // @[PPU.scala 53:26]
      scanlineY <= 9'h0; // @[PPU.scala 53:26]
    end else if (scanlineX == 9'h154) begin // @[PPU.scala 61:29]
      if (scanlineY == 9'h105) begin // @[PPU.scala 65:31]
        scanlineY <= 9'h0; // @[PPU.scala 66:17]
      end else begin
        scanlineY <= _scanlineY_T_1; // @[PPU.scala 63:15]
      end
    end
    if (reset) begin // @[PPU.scala 56:27]
      vblankFlag <= 1'h0; // @[PPU.scala 56:27]
    end else if (io_cpuRead) begin // @[PPU.scala 86:20]
      if (3'h2 == io_cpuAddr) begin // @[PPU.scala 87:24]
        vblankFlag <= 1'h0; // @[PPU.scala 90:20]
      end else begin
        vblankFlag <= _GEN_6;
      end
    end else begin
      vblankFlag <= _GEN_6;
    end
  end
endmodule
module MemoryController(
  input         clock,
  input  [15:0] io_cpuAddr,
  input  [7:0]  io_cpuDataIn,
  output [7:0]  io_cpuDataOut,
  input         io_cpuWrite,
  input         io_cpuRead,
  output [2:0]  io_ppuAddr,
  output [7:0]  io_ppuDataIn,
  input  [7:0]  io_ppuDataOut,
  output        io_ppuWrite,
  output        io_ppuRead,
  input  [7:0]  io_controller1,
  input  [7:0]  io_controller2
);
  reg [7:0] internalRAM [0:2047]; // @[MemoryController.scala 29:32]
  wire  internalRAM_io_cpuDataOut_MPORT_en; // @[MemoryController.scala 29:32]
  wire [10:0] internalRAM_io_cpuDataOut_MPORT_addr; // @[MemoryController.scala 29:32]
  wire [7:0] internalRAM_io_cpuDataOut_MPORT_data; // @[MemoryController.scala 29:32]
  wire [7:0] internalRAM_MPORT_data; // @[MemoryController.scala 29:32]
  wire [10:0] internalRAM_MPORT_addr; // @[MemoryController.scala 29:32]
  wire  internalRAM_MPORT_mask; // @[MemoryController.scala 29:32]
  wire  internalRAM_MPORT_en; // @[MemoryController.scala 29:32]
  reg  internalRAM_io_cpuDataOut_MPORT_en_pipe_0;
  reg [10:0] internalRAM_io_cpuDataOut_MPORT_addr_pipe_0;
  reg [7:0] prgROM [0:32767]; // @[MemoryController.scala 32:27]
  wire  prgROM_io_cpuDataOut_MPORT_1_en; // @[MemoryController.scala 32:27]
  wire [14:0] prgROM_io_cpuDataOut_MPORT_1_addr; // @[MemoryController.scala 32:27]
  wire [7:0] prgROM_io_cpuDataOut_MPORT_1_data; // @[MemoryController.scala 32:27]
  wire [7:0] prgROM_MPORT_1_data; // @[MemoryController.scala 32:27]
  wire [14:0] prgROM_MPORT_1_addr; // @[MemoryController.scala 32:27]
  wire  prgROM_MPORT_1_mask; // @[MemoryController.scala 32:27]
  wire  prgROM_MPORT_1_en; // @[MemoryController.scala 32:27]
  reg  prgROM_io_cpuDataOut_MPORT_1_en_pipe_0;
  reg [14:0] prgROM_io_cpuDataOut_MPORT_1_addr_pipe_0;
  wire  _T = io_cpuAddr < 16'h2000; // @[MemoryController.scala 51:21]
  wire  _T_3 = io_cpuAddr >= 16'h2000 & io_cpuAddr < 16'h4000; // @[MemoryController.scala 55:39]
  wire  _T_6 = io_cpuAddr >= 16'h8000; // @[MemoryController.scala 66:27]
  wire [15:0] romAddr = io_cpuAddr - 16'h8000; // @[MemoryController.scala 68:32]
  wire [7:0] _GEN_9 = io_cpuAddr >= 16'h8000 ? prgROM_io_cpuDataOut_MPORT_1_data : 8'h0; // @[MemoryController.scala 35:17 66:40 69:21]
  wire [7:0] _GEN_10 = io_cpuAddr == 16'h4017 ? io_controller2 : _GEN_9; // @[MemoryController.scala 63:41 65:21]
  wire  _GEN_11 = io_cpuAddr == 16'h4017 ? 1'h0 : _T_6; // @[MemoryController.scala 32:27 63:41]
  wire [7:0] _GEN_14 = io_cpuAddr == 16'h4016 ? io_controller1 : _GEN_10; // @[MemoryController.scala 60:41 62:21]
  wire  _GEN_15 = io_cpuAddr == 16'h4016 ? 1'h0 : _GEN_11; // @[MemoryController.scala 32:27 60:41]
  wire [2:0] _GEN_18 = io_cpuAddr >= 16'h2000 & io_cpuAddr < 16'h4000 ? io_cpuAddr[2:0] : 3'h0; // @[MemoryController.scala 36:14 55:65 57:18]
  wire [7:0] _GEN_20 = io_cpuAddr >= 16'h2000 & io_cpuAddr < 16'h4000 ? io_ppuDataOut : _GEN_14; // @[MemoryController.scala 55:65 59:21]
  wire  _GEN_21 = io_cpuAddr >= 16'h2000 & io_cpuAddr < 16'h4000 ? 1'h0 : _GEN_15; // @[MemoryController.scala 32:27 55:65]
  wire [7:0] _GEN_27 = io_cpuAddr < 16'h2000 ? internalRAM_io_cpuDataOut_MPORT_data : _GEN_20; // @[MemoryController.scala 51:33 54:21]
  wire [2:0] _GEN_28 = io_cpuAddr < 16'h2000 ? 3'h0 : _GEN_18; // @[MemoryController.scala 36:14 51:33]
  wire  _GEN_29 = io_cpuAddr < 16'h2000 ? 1'h0 : _T_3; // @[MemoryController.scala 39:14 51:33]
  wire  _GEN_30 = io_cpuAddr < 16'h2000 ? 1'h0 : _GEN_21; // @[MemoryController.scala 32:27 51:33]
  wire [2:0] _GEN_37 = io_cpuRead ? _GEN_28 : 3'h0; // @[MemoryController.scala 36:14 50:20]
  wire [2:0] _GEN_47 = _T_3 ? io_cpuAddr[2:0] : _GEN_37; // @[MemoryController.scala 78:65 80:18]
  wire [7:0] _GEN_48 = _T_3 ? io_cpuDataIn : 8'h0; // @[MemoryController.scala 37:16 78:65 81:20]
  wire  _GEN_52 = _T_3 ? 1'h0 : _T_6; // @[MemoryController.scala 32:27 78:65]
  wire [2:0] _GEN_60 = _T ? _GEN_37 : _GEN_47; // @[MemoryController.scala 74:33]
  wire [7:0] _GEN_61 = _T ? 8'h0 : _GEN_48; // @[MemoryController.scala 37:16 74:33]
  wire  _GEN_65 = _T ? 1'h0 : _GEN_52; // @[MemoryController.scala 32:27 74:33]
  assign internalRAM_io_cpuDataOut_MPORT_en = internalRAM_io_cpuDataOut_MPORT_en_pipe_0;
  assign internalRAM_io_cpuDataOut_MPORT_addr = internalRAM_io_cpuDataOut_MPORT_addr_pipe_0;
  assign internalRAM_io_cpuDataOut_MPORT_data = internalRAM[internalRAM_io_cpuDataOut_MPORT_addr]; // @[MemoryController.scala 29:32]
  assign internalRAM_MPORT_data = io_cpuDataIn;
  assign internalRAM_MPORT_addr = io_cpuAddr[10:0];
  assign internalRAM_MPORT_mask = 1'h1;
  assign internalRAM_MPORT_en = io_cpuWrite & _T;
  assign prgROM_io_cpuDataOut_MPORT_1_en = prgROM_io_cpuDataOut_MPORT_1_en_pipe_0;
  assign prgROM_io_cpuDataOut_MPORT_1_addr = prgROM_io_cpuDataOut_MPORT_1_addr_pipe_0;
  assign prgROM_io_cpuDataOut_MPORT_1_data = prgROM[prgROM_io_cpuDataOut_MPORT_1_addr]; // @[MemoryController.scala 32:27]
  assign prgROM_MPORT_1_data = io_cpuDataIn;
  assign prgROM_MPORT_1_addr = romAddr[14:0];
  assign prgROM_MPORT_1_mask = 1'h1;
  assign prgROM_MPORT_1_en = io_cpuWrite & _GEN_65;
  assign io_cpuDataOut = io_cpuRead ? _GEN_27 : 8'h0; // @[MemoryController.scala 35:17 50:20]
  assign io_ppuAddr = io_cpuWrite ? _GEN_60 : _GEN_37; // @[MemoryController.scala 73:21]
  assign io_ppuDataIn = io_cpuWrite ? _GEN_61 : 8'h0; // @[MemoryController.scala 37:16 73:21]
  assign io_ppuWrite = io_cpuWrite & _GEN_29; // @[MemoryController.scala 38:15 73:21]
  assign io_ppuRead = io_cpuRead & _GEN_29; // @[MemoryController.scala 39:14 50:20]
  always @(posedge clock) begin
    if (internalRAM_MPORT_en & internalRAM_MPORT_mask) begin
      internalRAM[internalRAM_MPORT_addr] <= internalRAM_MPORT_data; // @[MemoryController.scala 29:32]
    end
    internalRAM_io_cpuDataOut_MPORT_en_pipe_0 <= io_cpuRead & _T;
    if (io_cpuRead & _T) begin
      internalRAM_io_cpuDataOut_MPORT_addr_pipe_0 <= io_cpuAddr[10:0];
    end
    if (prgROM_MPORT_1_en & prgROM_MPORT_1_mask) begin
      prgROM[prgROM_MPORT_1_addr] <= prgROM_MPORT_1_data; // @[MemoryController.scala 32:27]
    end
    prgROM_io_cpuDataOut_MPORT_1_en_pipe_0 <= io_cpuRead & _GEN_30;
    if (io_cpuRead & _GEN_30) begin
      prgROM_io_cpuDataOut_MPORT_1_addr_pipe_0 <= romAddr[14:0];
    end
  end
endmodule
module NESSystem(
  input         clock,
  input         reset,
  output [8:0]  io_pixelX,
  output [8:0]  io_pixelY,
  output [5:0]  io_pixelColor,
  output        io_vblank,
  input  [7:0]  io_controller1,
  input  [7:0]  io_controller2,
  output [7:0]  io_debug_regA,
  output [7:0]  io_debug_regX,
  output [7:0]  io_debug_regY,
  output [15:0] io_debug_regPC,
  output [7:0]  io_debug_regSP,
  output        io_debug_flagC,
  output        io_debug_flagZ,
  output        io_debug_flagN,
  output        io_debug_flagV,
  output [7:0]  io_debug_opcode,
  input         io_romLoadEn,
  input  [15:0] io_romLoadAddr,
  input  [7:0]  io_romLoadData
);
  wire  cpu_clock; // @[NESSystem.scala 30:19]
  wire  cpu_reset; // @[NESSystem.scala 30:19]
  wire [15:0] cpu_io_memAddr; // @[NESSystem.scala 30:19]
  wire [7:0] cpu_io_memDataOut; // @[NESSystem.scala 30:19]
  wire [7:0] cpu_io_memDataIn; // @[NESSystem.scala 30:19]
  wire  cpu_io_memWrite; // @[NESSystem.scala 30:19]
  wire  cpu_io_memRead; // @[NESSystem.scala 30:19]
  wire [7:0] cpu_io_debug_regA; // @[NESSystem.scala 30:19]
  wire [7:0] cpu_io_debug_regX; // @[NESSystem.scala 30:19]
  wire [7:0] cpu_io_debug_regY; // @[NESSystem.scala 30:19]
  wire [15:0] cpu_io_debug_regPC; // @[NESSystem.scala 30:19]
  wire [7:0] cpu_io_debug_regSP; // @[NESSystem.scala 30:19]
  wire  cpu_io_debug_flagC; // @[NESSystem.scala 30:19]
  wire  cpu_io_debug_flagZ; // @[NESSystem.scala 30:19]
  wire  cpu_io_debug_flagN; // @[NESSystem.scala 30:19]
  wire  cpu_io_debug_flagV; // @[NESSystem.scala 30:19]
  wire [7:0] cpu_io_debug_opcode; // @[NESSystem.scala 30:19]
  wire  ppu_clock; // @[NESSystem.scala 31:19]
  wire  ppu_reset; // @[NESSystem.scala 31:19]
  wire [2:0] ppu_io_cpuAddr; // @[NESSystem.scala 31:19]
  wire [7:0] ppu_io_cpuDataIn; // @[NESSystem.scala 31:19]
  wire [7:0] ppu_io_cpuDataOut; // @[NESSystem.scala 31:19]
  wire  ppu_io_cpuWrite; // @[NESSystem.scala 31:19]
  wire  ppu_io_cpuRead; // @[NESSystem.scala 31:19]
  wire [8:0] ppu_io_pixelX; // @[NESSystem.scala 31:19]
  wire [8:0] ppu_io_pixelY; // @[NESSystem.scala 31:19]
  wire  ppu_io_vblank; // @[NESSystem.scala 31:19]
  wire  memory_clock; // @[NESSystem.scala 32:22]
  wire [15:0] memory_io_cpuAddr; // @[NESSystem.scala 32:22]
  wire [7:0] memory_io_cpuDataIn; // @[NESSystem.scala 32:22]
  wire [7:0] memory_io_cpuDataOut; // @[NESSystem.scala 32:22]
  wire  memory_io_cpuWrite; // @[NESSystem.scala 32:22]
  wire  memory_io_cpuRead; // @[NESSystem.scala 32:22]
  wire [2:0] memory_io_ppuAddr; // @[NESSystem.scala 32:22]
  wire [7:0] memory_io_ppuDataIn; // @[NESSystem.scala 32:22]
  wire [7:0] memory_io_ppuDataOut; // @[NESSystem.scala 32:22]
  wire  memory_io_ppuWrite; // @[NESSystem.scala 32:22]
  wire  memory_io_ppuRead; // @[NESSystem.scala 32:22]
  wire [7:0] memory_io_controller1; // @[NESSystem.scala 32:22]
  wire [7:0] memory_io_controller2; // @[NESSystem.scala 32:22]
  CPU6502 cpu ( // @[NESSystem.scala 30:19]
    .clock(cpu_clock),
    .reset(cpu_reset),
    .io_memAddr(cpu_io_memAddr),
    .io_memDataOut(cpu_io_memDataOut),
    .io_memDataIn(cpu_io_memDataIn),
    .io_memWrite(cpu_io_memWrite),
    .io_memRead(cpu_io_memRead),
    .io_debug_regA(cpu_io_debug_regA),
    .io_debug_regX(cpu_io_debug_regX),
    .io_debug_regY(cpu_io_debug_regY),
    .io_debug_regPC(cpu_io_debug_regPC),
    .io_debug_regSP(cpu_io_debug_regSP),
    .io_debug_flagC(cpu_io_debug_flagC),
    .io_debug_flagZ(cpu_io_debug_flagZ),
    .io_debug_flagN(cpu_io_debug_flagN),
    .io_debug_flagV(cpu_io_debug_flagV),
    .io_debug_opcode(cpu_io_debug_opcode)
  );
  PPU ppu ( // @[NESSystem.scala 31:19]
    .clock(ppu_clock),
    .reset(ppu_reset),
    .io_cpuAddr(ppu_io_cpuAddr),
    .io_cpuDataIn(ppu_io_cpuDataIn),
    .io_cpuDataOut(ppu_io_cpuDataOut),
    .io_cpuWrite(ppu_io_cpuWrite),
    .io_cpuRead(ppu_io_cpuRead),
    .io_pixelX(ppu_io_pixelX),
    .io_pixelY(ppu_io_pixelY),
    .io_vblank(ppu_io_vblank)
  );
  MemoryController memory ( // @[NESSystem.scala 32:22]
    .clock(memory_clock),
    .io_cpuAddr(memory_io_cpuAddr),
    .io_cpuDataIn(memory_io_cpuDataIn),
    .io_cpuDataOut(memory_io_cpuDataOut),
    .io_cpuWrite(memory_io_cpuWrite),
    .io_cpuRead(memory_io_cpuRead),
    .io_ppuAddr(memory_io_ppuAddr),
    .io_ppuDataIn(memory_io_ppuDataIn),
    .io_ppuDataOut(memory_io_ppuDataOut),
    .io_ppuWrite(memory_io_ppuWrite),
    .io_ppuRead(memory_io_ppuRead),
    .io_controller1(memory_io_controller1),
    .io_controller2(memory_io_controller2)
  );
  assign io_pixelX = ppu_io_pixelX; // @[NESSystem.scala 53:13]
  assign io_pixelY = ppu_io_pixelY; // @[NESSystem.scala 54:13]
  assign io_pixelColor = 6'h0; // @[NESSystem.scala 55:17]
  assign io_vblank = ppu_io_vblank; // @[NESSystem.scala 56:13]
  assign io_debug_regA = cpu_io_debug_regA; // @[NESSystem.scala 59:12]
  assign io_debug_regX = cpu_io_debug_regX; // @[NESSystem.scala 59:12]
  assign io_debug_regY = cpu_io_debug_regY; // @[NESSystem.scala 59:12]
  assign io_debug_regPC = cpu_io_debug_regPC; // @[NESSystem.scala 59:12]
  assign io_debug_regSP = cpu_io_debug_regSP; // @[NESSystem.scala 59:12]
  assign io_debug_flagC = cpu_io_debug_flagC; // @[NESSystem.scala 59:12]
  assign io_debug_flagZ = cpu_io_debug_flagZ; // @[NESSystem.scala 59:12]
  assign io_debug_flagN = cpu_io_debug_flagN; // @[NESSystem.scala 59:12]
  assign io_debug_flagV = cpu_io_debug_flagV; // @[NESSystem.scala 59:12]
  assign io_debug_opcode = cpu_io_debug_opcode; // @[NESSystem.scala 59:12]
  assign cpu_clock = clock;
  assign cpu_reset = reset;
  assign cpu_io_memDataIn = memory_io_cpuDataOut; // @[NESSystem.scala 37:20]
  assign ppu_clock = clock;
  assign ppu_reset = reset;
  assign ppu_io_cpuAddr = memory_io_ppuAddr; // @[NESSystem.scala 42:18]
  assign ppu_io_cpuDataIn = memory_io_ppuDataIn; // @[NESSystem.scala 43:20]
  assign ppu_io_cpuWrite = memory_io_ppuWrite; // @[NESSystem.scala 45:19]
  assign ppu_io_cpuRead = memory_io_ppuRead; // @[NESSystem.scala 46:18]
  assign memory_clock = clock;
  assign memory_io_cpuAddr = cpu_io_memAddr; // @[NESSystem.scala 35:21]
  assign memory_io_cpuDataIn = cpu_io_memDataOut; // @[NESSystem.scala 36:23]
  assign memory_io_cpuWrite = cpu_io_memWrite; // @[NESSystem.scala 38:22]
  assign memory_io_cpuRead = cpu_io_memRead; // @[NESSystem.scala 39:21]
  assign memory_io_ppuDataOut = ppu_io_cpuDataOut; // @[NESSystem.scala 44:24]
  assign memory_io_controller1 = io_controller1; // @[NESSystem.scala 49:25]
  assign memory_io_controller2 = io_controller2; // @[NESSystem.scala 50:25]
endmodule
